magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< metal3 >>
rect -2550 2472 2549 2500
rect -2550 2408 2465 2472
rect 2529 2408 2549 2472
rect -2550 2392 2549 2408
rect -2550 2328 2465 2392
rect 2529 2328 2549 2392
rect -2550 2312 2549 2328
rect -2550 2248 2465 2312
rect 2529 2248 2549 2312
rect -2550 2232 2549 2248
rect -2550 2168 2465 2232
rect 2529 2168 2549 2232
rect -2550 2152 2549 2168
rect -2550 2088 2465 2152
rect 2529 2088 2549 2152
rect -2550 2072 2549 2088
rect -2550 2008 2465 2072
rect 2529 2008 2549 2072
rect -2550 1992 2549 2008
rect -2550 1928 2465 1992
rect 2529 1928 2549 1992
rect -2550 1912 2549 1928
rect -2550 1848 2465 1912
rect 2529 1848 2549 1912
rect -2550 1832 2549 1848
rect -2550 1768 2465 1832
rect 2529 1768 2549 1832
rect -2550 1752 2549 1768
rect -2550 1688 2465 1752
rect 2529 1688 2549 1752
rect -2550 1672 2549 1688
rect -2550 1608 2465 1672
rect 2529 1608 2549 1672
rect -2550 1592 2549 1608
rect -2550 1528 2465 1592
rect 2529 1528 2549 1592
rect -2550 1512 2549 1528
rect -2550 1448 2465 1512
rect 2529 1448 2549 1512
rect -2550 1432 2549 1448
rect -2550 1368 2465 1432
rect 2529 1368 2549 1432
rect -2550 1352 2549 1368
rect -2550 1288 2465 1352
rect 2529 1288 2549 1352
rect -2550 1272 2549 1288
rect -2550 1208 2465 1272
rect 2529 1208 2549 1272
rect -2550 1192 2549 1208
rect -2550 1128 2465 1192
rect 2529 1128 2549 1192
rect -2550 1112 2549 1128
rect -2550 1048 2465 1112
rect 2529 1048 2549 1112
rect -2550 1032 2549 1048
rect -2550 968 2465 1032
rect 2529 968 2549 1032
rect -2550 952 2549 968
rect -2550 888 2465 952
rect 2529 888 2549 952
rect -2550 872 2549 888
rect -2550 808 2465 872
rect 2529 808 2549 872
rect -2550 792 2549 808
rect -2550 728 2465 792
rect 2529 728 2549 792
rect -2550 712 2549 728
rect -2550 648 2465 712
rect 2529 648 2549 712
rect -2550 632 2549 648
rect -2550 568 2465 632
rect 2529 568 2549 632
rect -2550 552 2549 568
rect -2550 488 2465 552
rect 2529 488 2549 552
rect -2550 472 2549 488
rect -2550 408 2465 472
rect 2529 408 2549 472
rect -2550 392 2549 408
rect -2550 328 2465 392
rect 2529 328 2549 392
rect -2550 312 2549 328
rect -2550 248 2465 312
rect 2529 248 2549 312
rect -2550 232 2549 248
rect -2550 168 2465 232
rect 2529 168 2549 232
rect -2550 152 2549 168
rect -2550 88 2465 152
rect 2529 88 2549 152
rect -2550 72 2549 88
rect -2550 8 2465 72
rect 2529 8 2549 72
rect -2550 -8 2549 8
rect -2550 -72 2465 -8
rect 2529 -72 2549 -8
rect -2550 -88 2549 -72
rect -2550 -152 2465 -88
rect 2529 -152 2549 -88
rect -2550 -168 2549 -152
rect -2550 -232 2465 -168
rect 2529 -232 2549 -168
rect -2550 -248 2549 -232
rect -2550 -312 2465 -248
rect 2529 -312 2549 -248
rect -2550 -328 2549 -312
rect -2550 -392 2465 -328
rect 2529 -392 2549 -328
rect -2550 -408 2549 -392
rect -2550 -472 2465 -408
rect 2529 -472 2549 -408
rect -2550 -488 2549 -472
rect -2550 -552 2465 -488
rect 2529 -552 2549 -488
rect -2550 -568 2549 -552
rect -2550 -632 2465 -568
rect 2529 -632 2549 -568
rect -2550 -648 2549 -632
rect -2550 -712 2465 -648
rect 2529 -712 2549 -648
rect -2550 -728 2549 -712
rect -2550 -792 2465 -728
rect 2529 -792 2549 -728
rect -2550 -808 2549 -792
rect -2550 -872 2465 -808
rect 2529 -872 2549 -808
rect -2550 -888 2549 -872
rect -2550 -952 2465 -888
rect 2529 -952 2549 -888
rect -2550 -968 2549 -952
rect -2550 -1032 2465 -968
rect 2529 -1032 2549 -968
rect -2550 -1048 2549 -1032
rect -2550 -1112 2465 -1048
rect 2529 -1112 2549 -1048
rect -2550 -1128 2549 -1112
rect -2550 -1192 2465 -1128
rect 2529 -1192 2549 -1128
rect -2550 -1208 2549 -1192
rect -2550 -1272 2465 -1208
rect 2529 -1272 2549 -1208
rect -2550 -1288 2549 -1272
rect -2550 -1352 2465 -1288
rect 2529 -1352 2549 -1288
rect -2550 -1368 2549 -1352
rect -2550 -1432 2465 -1368
rect 2529 -1432 2549 -1368
rect -2550 -1448 2549 -1432
rect -2550 -1512 2465 -1448
rect 2529 -1512 2549 -1448
rect -2550 -1528 2549 -1512
rect -2550 -1592 2465 -1528
rect 2529 -1592 2549 -1528
rect -2550 -1608 2549 -1592
rect -2550 -1672 2465 -1608
rect 2529 -1672 2549 -1608
rect -2550 -1688 2549 -1672
rect -2550 -1752 2465 -1688
rect 2529 -1752 2549 -1688
rect -2550 -1768 2549 -1752
rect -2550 -1832 2465 -1768
rect 2529 -1832 2549 -1768
rect -2550 -1848 2549 -1832
rect -2550 -1912 2465 -1848
rect 2529 -1912 2549 -1848
rect -2550 -1928 2549 -1912
rect -2550 -1992 2465 -1928
rect 2529 -1992 2549 -1928
rect -2550 -2008 2549 -1992
rect -2550 -2072 2465 -2008
rect 2529 -2072 2549 -2008
rect -2550 -2088 2549 -2072
rect -2550 -2152 2465 -2088
rect 2529 -2152 2549 -2088
rect -2550 -2168 2549 -2152
rect -2550 -2232 2465 -2168
rect 2529 -2232 2549 -2168
rect -2550 -2248 2549 -2232
rect -2550 -2312 2465 -2248
rect 2529 -2312 2549 -2248
rect -2550 -2328 2549 -2312
rect -2550 -2392 2465 -2328
rect 2529 -2392 2549 -2328
rect -2550 -2408 2549 -2392
rect -2550 -2472 2465 -2408
rect 2529 -2472 2549 -2408
rect -2550 -2500 2549 -2472
<< via3 >>
rect 2465 2408 2529 2472
rect 2465 2328 2529 2392
rect 2465 2248 2529 2312
rect 2465 2168 2529 2232
rect 2465 2088 2529 2152
rect 2465 2008 2529 2072
rect 2465 1928 2529 1992
rect 2465 1848 2529 1912
rect 2465 1768 2529 1832
rect 2465 1688 2529 1752
rect 2465 1608 2529 1672
rect 2465 1528 2529 1592
rect 2465 1448 2529 1512
rect 2465 1368 2529 1432
rect 2465 1288 2529 1352
rect 2465 1208 2529 1272
rect 2465 1128 2529 1192
rect 2465 1048 2529 1112
rect 2465 968 2529 1032
rect 2465 888 2529 952
rect 2465 808 2529 872
rect 2465 728 2529 792
rect 2465 648 2529 712
rect 2465 568 2529 632
rect 2465 488 2529 552
rect 2465 408 2529 472
rect 2465 328 2529 392
rect 2465 248 2529 312
rect 2465 168 2529 232
rect 2465 88 2529 152
rect 2465 8 2529 72
rect 2465 -72 2529 -8
rect 2465 -152 2529 -88
rect 2465 -232 2529 -168
rect 2465 -312 2529 -248
rect 2465 -392 2529 -328
rect 2465 -472 2529 -408
rect 2465 -552 2529 -488
rect 2465 -632 2529 -568
rect 2465 -712 2529 -648
rect 2465 -792 2529 -728
rect 2465 -872 2529 -808
rect 2465 -952 2529 -888
rect 2465 -1032 2529 -968
rect 2465 -1112 2529 -1048
rect 2465 -1192 2529 -1128
rect 2465 -1272 2529 -1208
rect 2465 -1352 2529 -1288
rect 2465 -1432 2529 -1368
rect 2465 -1512 2529 -1448
rect 2465 -1592 2529 -1528
rect 2465 -1672 2529 -1608
rect 2465 -1752 2529 -1688
rect 2465 -1832 2529 -1768
rect 2465 -1912 2529 -1848
rect 2465 -1992 2529 -1928
rect 2465 -2072 2529 -2008
rect 2465 -2152 2529 -2088
rect 2465 -2232 2529 -2168
rect 2465 -2312 2529 -2248
rect 2465 -2392 2529 -2328
rect 2465 -2472 2529 -2408
<< mimcap >>
rect -2450 2352 2350 2400
rect -2450 -2352 -2402 2352
rect 2302 -2352 2350 2352
rect -2450 -2400 2350 -2352
<< mimcapcontact >>
rect -2402 -2352 2302 2352
<< metal4 >>
rect 2449 2472 2545 2488
rect 2449 2408 2465 2472
rect 2529 2408 2545 2472
rect 2449 2392 2545 2408
rect -2411 2352 2311 2361
rect -2411 -2352 -2402 2352
rect 2302 -2352 2311 2352
rect -2411 -2361 2311 -2352
rect 2449 2328 2465 2392
rect 2529 2328 2545 2392
rect 2449 2312 2545 2328
rect 2449 2248 2465 2312
rect 2529 2248 2545 2312
rect 2449 2232 2545 2248
rect 2449 2168 2465 2232
rect 2529 2168 2545 2232
rect 2449 2152 2545 2168
rect 2449 2088 2465 2152
rect 2529 2088 2545 2152
rect 2449 2072 2545 2088
rect 2449 2008 2465 2072
rect 2529 2008 2545 2072
rect 2449 1992 2545 2008
rect 2449 1928 2465 1992
rect 2529 1928 2545 1992
rect 2449 1912 2545 1928
rect 2449 1848 2465 1912
rect 2529 1848 2545 1912
rect 2449 1832 2545 1848
rect 2449 1768 2465 1832
rect 2529 1768 2545 1832
rect 2449 1752 2545 1768
rect 2449 1688 2465 1752
rect 2529 1688 2545 1752
rect 2449 1672 2545 1688
rect 2449 1608 2465 1672
rect 2529 1608 2545 1672
rect 2449 1592 2545 1608
rect 2449 1528 2465 1592
rect 2529 1528 2545 1592
rect 2449 1512 2545 1528
rect 2449 1448 2465 1512
rect 2529 1448 2545 1512
rect 2449 1432 2545 1448
rect 2449 1368 2465 1432
rect 2529 1368 2545 1432
rect 2449 1352 2545 1368
rect 2449 1288 2465 1352
rect 2529 1288 2545 1352
rect 2449 1272 2545 1288
rect 2449 1208 2465 1272
rect 2529 1208 2545 1272
rect 2449 1192 2545 1208
rect 2449 1128 2465 1192
rect 2529 1128 2545 1192
rect 2449 1112 2545 1128
rect 2449 1048 2465 1112
rect 2529 1048 2545 1112
rect 2449 1032 2545 1048
rect 2449 968 2465 1032
rect 2529 968 2545 1032
rect 2449 952 2545 968
rect 2449 888 2465 952
rect 2529 888 2545 952
rect 2449 872 2545 888
rect 2449 808 2465 872
rect 2529 808 2545 872
rect 2449 792 2545 808
rect 2449 728 2465 792
rect 2529 728 2545 792
rect 2449 712 2545 728
rect 2449 648 2465 712
rect 2529 648 2545 712
rect 2449 632 2545 648
rect 2449 568 2465 632
rect 2529 568 2545 632
rect 2449 552 2545 568
rect 2449 488 2465 552
rect 2529 488 2545 552
rect 2449 472 2545 488
rect 2449 408 2465 472
rect 2529 408 2545 472
rect 2449 392 2545 408
rect 2449 328 2465 392
rect 2529 328 2545 392
rect 2449 312 2545 328
rect 2449 248 2465 312
rect 2529 248 2545 312
rect 2449 232 2545 248
rect 2449 168 2465 232
rect 2529 168 2545 232
rect 2449 152 2545 168
rect 2449 88 2465 152
rect 2529 88 2545 152
rect 2449 72 2545 88
rect 2449 8 2465 72
rect 2529 8 2545 72
rect 2449 -8 2545 8
rect 2449 -72 2465 -8
rect 2529 -72 2545 -8
rect 2449 -88 2545 -72
rect 2449 -152 2465 -88
rect 2529 -152 2545 -88
rect 2449 -168 2545 -152
rect 2449 -232 2465 -168
rect 2529 -232 2545 -168
rect 2449 -248 2545 -232
rect 2449 -312 2465 -248
rect 2529 -312 2545 -248
rect 2449 -328 2545 -312
rect 2449 -392 2465 -328
rect 2529 -392 2545 -328
rect 2449 -408 2545 -392
rect 2449 -472 2465 -408
rect 2529 -472 2545 -408
rect 2449 -488 2545 -472
rect 2449 -552 2465 -488
rect 2529 -552 2545 -488
rect 2449 -568 2545 -552
rect 2449 -632 2465 -568
rect 2529 -632 2545 -568
rect 2449 -648 2545 -632
rect 2449 -712 2465 -648
rect 2529 -712 2545 -648
rect 2449 -728 2545 -712
rect 2449 -792 2465 -728
rect 2529 -792 2545 -728
rect 2449 -808 2545 -792
rect 2449 -872 2465 -808
rect 2529 -872 2545 -808
rect 2449 -888 2545 -872
rect 2449 -952 2465 -888
rect 2529 -952 2545 -888
rect 2449 -968 2545 -952
rect 2449 -1032 2465 -968
rect 2529 -1032 2545 -968
rect 2449 -1048 2545 -1032
rect 2449 -1112 2465 -1048
rect 2529 -1112 2545 -1048
rect 2449 -1128 2545 -1112
rect 2449 -1192 2465 -1128
rect 2529 -1192 2545 -1128
rect 2449 -1208 2545 -1192
rect 2449 -1272 2465 -1208
rect 2529 -1272 2545 -1208
rect 2449 -1288 2545 -1272
rect 2449 -1352 2465 -1288
rect 2529 -1352 2545 -1288
rect 2449 -1368 2545 -1352
rect 2449 -1432 2465 -1368
rect 2529 -1432 2545 -1368
rect 2449 -1448 2545 -1432
rect 2449 -1512 2465 -1448
rect 2529 -1512 2545 -1448
rect 2449 -1528 2545 -1512
rect 2449 -1592 2465 -1528
rect 2529 -1592 2545 -1528
rect 2449 -1608 2545 -1592
rect 2449 -1672 2465 -1608
rect 2529 -1672 2545 -1608
rect 2449 -1688 2545 -1672
rect 2449 -1752 2465 -1688
rect 2529 -1752 2545 -1688
rect 2449 -1768 2545 -1752
rect 2449 -1832 2465 -1768
rect 2529 -1832 2545 -1768
rect 2449 -1848 2545 -1832
rect 2449 -1912 2465 -1848
rect 2529 -1912 2545 -1848
rect 2449 -1928 2545 -1912
rect 2449 -1992 2465 -1928
rect 2529 -1992 2545 -1928
rect 2449 -2008 2545 -1992
rect 2449 -2072 2465 -2008
rect 2529 -2072 2545 -2008
rect 2449 -2088 2545 -2072
rect 2449 -2152 2465 -2088
rect 2529 -2152 2545 -2088
rect 2449 -2168 2545 -2152
rect 2449 -2232 2465 -2168
rect 2529 -2232 2545 -2168
rect 2449 -2248 2545 -2232
rect 2449 -2312 2465 -2248
rect 2529 -2312 2545 -2248
rect 2449 -2328 2545 -2312
rect 2449 -2392 2465 -2328
rect 2529 -2392 2545 -2328
rect 2449 -2408 2545 -2392
rect 2449 -2472 2465 -2408
rect 2529 -2472 2545 -2408
rect 2449 -2488 2545 -2472
<< properties >>
string FIXED_BBOX -2550 -2500 2450 2500
<< end >>
