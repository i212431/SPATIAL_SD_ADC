magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< metal3 >>
rect -1650 1552 1649 1600
rect -1650 1488 1565 1552
rect 1629 1488 1649 1552
rect -1650 1472 1649 1488
rect -1650 1408 1565 1472
rect 1629 1408 1649 1472
rect -1650 1392 1649 1408
rect -1650 1328 1565 1392
rect 1629 1328 1649 1392
rect -1650 1312 1649 1328
rect -1650 1248 1565 1312
rect 1629 1248 1649 1312
rect -1650 1232 1649 1248
rect -1650 1168 1565 1232
rect 1629 1168 1649 1232
rect -1650 1152 1649 1168
rect -1650 1088 1565 1152
rect 1629 1088 1649 1152
rect -1650 1072 1649 1088
rect -1650 1008 1565 1072
rect 1629 1008 1649 1072
rect -1650 992 1649 1008
rect -1650 928 1565 992
rect 1629 928 1649 992
rect -1650 912 1649 928
rect -1650 848 1565 912
rect 1629 848 1649 912
rect -1650 832 1649 848
rect -1650 768 1565 832
rect 1629 768 1649 832
rect -1650 752 1649 768
rect -1650 688 1565 752
rect 1629 688 1649 752
rect -1650 672 1649 688
rect -1650 608 1565 672
rect 1629 608 1649 672
rect -1650 592 1649 608
rect -1650 528 1565 592
rect 1629 528 1649 592
rect -1650 512 1649 528
rect -1650 448 1565 512
rect 1629 448 1649 512
rect -1650 432 1649 448
rect -1650 368 1565 432
rect 1629 368 1649 432
rect -1650 352 1649 368
rect -1650 288 1565 352
rect 1629 288 1649 352
rect -1650 272 1649 288
rect -1650 208 1565 272
rect 1629 208 1649 272
rect -1650 192 1649 208
rect -1650 128 1565 192
rect 1629 128 1649 192
rect -1650 112 1649 128
rect -1650 48 1565 112
rect 1629 48 1649 112
rect -1650 32 1649 48
rect -1650 -32 1565 32
rect 1629 -32 1649 32
rect -1650 -48 1649 -32
rect -1650 -112 1565 -48
rect 1629 -112 1649 -48
rect -1650 -128 1649 -112
rect -1650 -192 1565 -128
rect 1629 -192 1649 -128
rect -1650 -208 1649 -192
rect -1650 -272 1565 -208
rect 1629 -272 1649 -208
rect -1650 -288 1649 -272
rect -1650 -352 1565 -288
rect 1629 -352 1649 -288
rect -1650 -368 1649 -352
rect -1650 -432 1565 -368
rect 1629 -432 1649 -368
rect -1650 -448 1649 -432
rect -1650 -512 1565 -448
rect 1629 -512 1649 -448
rect -1650 -528 1649 -512
rect -1650 -592 1565 -528
rect 1629 -592 1649 -528
rect -1650 -608 1649 -592
rect -1650 -672 1565 -608
rect 1629 -672 1649 -608
rect -1650 -688 1649 -672
rect -1650 -752 1565 -688
rect 1629 -752 1649 -688
rect -1650 -768 1649 -752
rect -1650 -832 1565 -768
rect 1629 -832 1649 -768
rect -1650 -848 1649 -832
rect -1650 -912 1565 -848
rect 1629 -912 1649 -848
rect -1650 -928 1649 -912
rect -1650 -992 1565 -928
rect 1629 -992 1649 -928
rect -1650 -1008 1649 -992
rect -1650 -1072 1565 -1008
rect 1629 -1072 1649 -1008
rect -1650 -1088 1649 -1072
rect -1650 -1152 1565 -1088
rect 1629 -1152 1649 -1088
rect -1650 -1168 1649 -1152
rect -1650 -1232 1565 -1168
rect 1629 -1232 1649 -1168
rect -1650 -1248 1649 -1232
rect -1650 -1312 1565 -1248
rect 1629 -1312 1649 -1248
rect -1650 -1328 1649 -1312
rect -1650 -1392 1565 -1328
rect 1629 -1392 1649 -1328
rect -1650 -1408 1649 -1392
rect -1650 -1472 1565 -1408
rect 1629 -1472 1649 -1408
rect -1650 -1488 1649 -1472
rect -1650 -1552 1565 -1488
rect 1629 -1552 1649 -1488
rect -1650 -1600 1649 -1552
<< via3 >>
rect 1565 1488 1629 1552
rect 1565 1408 1629 1472
rect 1565 1328 1629 1392
rect 1565 1248 1629 1312
rect 1565 1168 1629 1232
rect 1565 1088 1629 1152
rect 1565 1008 1629 1072
rect 1565 928 1629 992
rect 1565 848 1629 912
rect 1565 768 1629 832
rect 1565 688 1629 752
rect 1565 608 1629 672
rect 1565 528 1629 592
rect 1565 448 1629 512
rect 1565 368 1629 432
rect 1565 288 1629 352
rect 1565 208 1629 272
rect 1565 128 1629 192
rect 1565 48 1629 112
rect 1565 -32 1629 32
rect 1565 -112 1629 -48
rect 1565 -192 1629 -128
rect 1565 -272 1629 -208
rect 1565 -352 1629 -288
rect 1565 -432 1629 -368
rect 1565 -512 1629 -448
rect 1565 -592 1629 -528
rect 1565 -672 1629 -608
rect 1565 -752 1629 -688
rect 1565 -832 1629 -768
rect 1565 -912 1629 -848
rect 1565 -992 1629 -928
rect 1565 -1072 1629 -1008
rect 1565 -1152 1629 -1088
rect 1565 -1232 1629 -1168
rect 1565 -1312 1629 -1248
rect 1565 -1392 1629 -1328
rect 1565 -1472 1629 -1408
rect 1565 -1552 1629 -1488
<< mimcap >>
rect -1550 1432 1450 1500
rect -1550 -1432 -1482 1432
rect 1382 -1432 1450 1432
rect -1550 -1500 1450 -1432
<< mimcapcontact >>
rect -1482 -1432 1382 1432
<< metal4 >>
rect 1549 1552 1645 1588
rect 1549 1488 1565 1552
rect 1629 1488 1645 1552
rect 1549 1472 1645 1488
rect -1511 1432 1411 1461
rect -1511 -1432 -1482 1432
rect 1382 -1432 1411 1432
rect -1511 -1461 1411 -1432
rect 1549 1408 1565 1472
rect 1629 1408 1645 1472
rect 1549 1392 1645 1408
rect 1549 1328 1565 1392
rect 1629 1328 1645 1392
rect 1549 1312 1645 1328
rect 1549 1248 1565 1312
rect 1629 1248 1645 1312
rect 1549 1232 1645 1248
rect 1549 1168 1565 1232
rect 1629 1168 1645 1232
rect 1549 1152 1645 1168
rect 1549 1088 1565 1152
rect 1629 1088 1645 1152
rect 1549 1072 1645 1088
rect 1549 1008 1565 1072
rect 1629 1008 1645 1072
rect 1549 992 1645 1008
rect 1549 928 1565 992
rect 1629 928 1645 992
rect 1549 912 1645 928
rect 1549 848 1565 912
rect 1629 848 1645 912
rect 1549 832 1645 848
rect 1549 768 1565 832
rect 1629 768 1645 832
rect 1549 752 1645 768
rect 1549 688 1565 752
rect 1629 688 1645 752
rect 1549 672 1645 688
rect 1549 608 1565 672
rect 1629 608 1645 672
rect 1549 592 1645 608
rect 1549 528 1565 592
rect 1629 528 1645 592
rect 1549 512 1645 528
rect 1549 448 1565 512
rect 1629 448 1645 512
rect 1549 432 1645 448
rect 1549 368 1565 432
rect 1629 368 1645 432
rect 1549 352 1645 368
rect 1549 288 1565 352
rect 1629 288 1645 352
rect 1549 272 1645 288
rect 1549 208 1565 272
rect 1629 208 1645 272
rect 1549 192 1645 208
rect 1549 128 1565 192
rect 1629 128 1645 192
rect 1549 112 1645 128
rect 1549 48 1565 112
rect 1629 48 1645 112
rect 1549 32 1645 48
rect 1549 -32 1565 32
rect 1629 -32 1645 32
rect 1549 -48 1645 -32
rect 1549 -112 1565 -48
rect 1629 -112 1645 -48
rect 1549 -128 1645 -112
rect 1549 -192 1565 -128
rect 1629 -192 1645 -128
rect 1549 -208 1645 -192
rect 1549 -272 1565 -208
rect 1629 -272 1645 -208
rect 1549 -288 1645 -272
rect 1549 -352 1565 -288
rect 1629 -352 1645 -288
rect 1549 -368 1645 -352
rect 1549 -432 1565 -368
rect 1629 -432 1645 -368
rect 1549 -448 1645 -432
rect 1549 -512 1565 -448
rect 1629 -512 1645 -448
rect 1549 -528 1645 -512
rect 1549 -592 1565 -528
rect 1629 -592 1645 -528
rect 1549 -608 1645 -592
rect 1549 -672 1565 -608
rect 1629 -672 1645 -608
rect 1549 -688 1645 -672
rect 1549 -752 1565 -688
rect 1629 -752 1645 -688
rect 1549 -768 1645 -752
rect 1549 -832 1565 -768
rect 1629 -832 1645 -768
rect 1549 -848 1645 -832
rect 1549 -912 1565 -848
rect 1629 -912 1645 -848
rect 1549 -928 1645 -912
rect 1549 -992 1565 -928
rect 1629 -992 1645 -928
rect 1549 -1008 1645 -992
rect 1549 -1072 1565 -1008
rect 1629 -1072 1645 -1008
rect 1549 -1088 1645 -1072
rect 1549 -1152 1565 -1088
rect 1629 -1152 1645 -1088
rect 1549 -1168 1645 -1152
rect 1549 -1232 1565 -1168
rect 1629 -1232 1645 -1168
rect 1549 -1248 1645 -1232
rect 1549 -1312 1565 -1248
rect 1629 -1312 1645 -1248
rect 1549 -1328 1645 -1312
rect 1549 -1392 1565 -1328
rect 1629 -1392 1645 -1328
rect 1549 -1408 1645 -1392
rect 1549 -1472 1565 -1408
rect 1629 -1472 1645 -1408
rect 1549 -1488 1645 -1472
rect 1549 -1552 1565 -1488
rect 1629 -1552 1645 -1488
rect 1549 -1588 1645 -1552
<< properties >>
string FIXED_BBOX -1650 -1600 1550 1600
<< end >>
