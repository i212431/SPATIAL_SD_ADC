magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< metal3 >>
rect -3150 1072 3149 1100
rect -3150 1008 3065 1072
rect 3129 1008 3149 1072
rect -3150 992 3149 1008
rect -3150 928 3065 992
rect 3129 928 3149 992
rect -3150 912 3149 928
rect -3150 848 3065 912
rect 3129 848 3149 912
rect -3150 832 3149 848
rect -3150 768 3065 832
rect 3129 768 3149 832
rect -3150 752 3149 768
rect -3150 688 3065 752
rect 3129 688 3149 752
rect -3150 672 3149 688
rect -3150 608 3065 672
rect 3129 608 3149 672
rect -3150 592 3149 608
rect -3150 528 3065 592
rect 3129 528 3149 592
rect -3150 512 3149 528
rect -3150 448 3065 512
rect 3129 448 3149 512
rect -3150 432 3149 448
rect -3150 368 3065 432
rect 3129 368 3149 432
rect -3150 352 3149 368
rect -3150 288 3065 352
rect 3129 288 3149 352
rect -3150 272 3149 288
rect -3150 208 3065 272
rect 3129 208 3149 272
rect -3150 192 3149 208
rect -3150 128 3065 192
rect 3129 128 3149 192
rect -3150 112 3149 128
rect -3150 48 3065 112
rect 3129 48 3149 112
rect -3150 32 3149 48
rect -3150 -32 3065 32
rect 3129 -32 3149 32
rect -3150 -48 3149 -32
rect -3150 -112 3065 -48
rect 3129 -112 3149 -48
rect -3150 -128 3149 -112
rect -3150 -192 3065 -128
rect 3129 -192 3149 -128
rect -3150 -208 3149 -192
rect -3150 -272 3065 -208
rect 3129 -272 3149 -208
rect -3150 -288 3149 -272
rect -3150 -352 3065 -288
rect 3129 -352 3149 -288
rect -3150 -368 3149 -352
rect -3150 -432 3065 -368
rect 3129 -432 3149 -368
rect -3150 -448 3149 -432
rect -3150 -512 3065 -448
rect 3129 -512 3149 -448
rect -3150 -528 3149 -512
rect -3150 -592 3065 -528
rect 3129 -592 3149 -528
rect -3150 -608 3149 -592
rect -3150 -672 3065 -608
rect 3129 -672 3149 -608
rect -3150 -688 3149 -672
rect -3150 -752 3065 -688
rect 3129 -752 3149 -688
rect -3150 -768 3149 -752
rect -3150 -832 3065 -768
rect 3129 -832 3149 -768
rect -3150 -848 3149 -832
rect -3150 -912 3065 -848
rect 3129 -912 3149 -848
rect -3150 -928 3149 -912
rect -3150 -992 3065 -928
rect 3129 -992 3149 -928
rect -3150 -1008 3149 -992
rect -3150 -1072 3065 -1008
rect 3129 -1072 3149 -1008
rect -3150 -1100 3149 -1072
<< via3 >>
rect 3065 1008 3129 1072
rect 3065 928 3129 992
rect 3065 848 3129 912
rect 3065 768 3129 832
rect 3065 688 3129 752
rect 3065 608 3129 672
rect 3065 528 3129 592
rect 3065 448 3129 512
rect 3065 368 3129 432
rect 3065 288 3129 352
rect 3065 208 3129 272
rect 3065 128 3129 192
rect 3065 48 3129 112
rect 3065 -32 3129 32
rect 3065 -112 3129 -48
rect 3065 -192 3129 -128
rect 3065 -272 3129 -208
rect 3065 -352 3129 -288
rect 3065 -432 3129 -368
rect 3065 -512 3129 -448
rect 3065 -592 3129 -528
rect 3065 -672 3129 -608
rect 3065 -752 3129 -688
rect 3065 -832 3129 -768
rect 3065 -912 3129 -848
rect 3065 -992 3129 -928
rect 3065 -1072 3129 -1008
<< mimcap >>
rect -3050 952 2950 1000
rect -3050 -952 -3002 952
rect 2902 -952 2950 952
rect -3050 -1000 2950 -952
<< mimcapcontact >>
rect -3002 -952 2902 952
<< metal4 >>
rect 3049 1072 3145 1088
rect 3049 1008 3065 1072
rect 3129 1008 3145 1072
rect 3049 992 3145 1008
rect -3011 952 2911 961
rect -3011 -952 -3002 952
rect 2902 -952 2911 952
rect -3011 -961 2911 -952
rect 3049 928 3065 992
rect 3129 928 3145 992
rect 3049 912 3145 928
rect 3049 848 3065 912
rect 3129 848 3145 912
rect 3049 832 3145 848
rect 3049 768 3065 832
rect 3129 768 3145 832
rect 3049 752 3145 768
rect 3049 688 3065 752
rect 3129 688 3145 752
rect 3049 672 3145 688
rect 3049 608 3065 672
rect 3129 608 3145 672
rect 3049 592 3145 608
rect 3049 528 3065 592
rect 3129 528 3145 592
rect 3049 512 3145 528
rect 3049 448 3065 512
rect 3129 448 3145 512
rect 3049 432 3145 448
rect 3049 368 3065 432
rect 3129 368 3145 432
rect 3049 352 3145 368
rect 3049 288 3065 352
rect 3129 288 3145 352
rect 3049 272 3145 288
rect 3049 208 3065 272
rect 3129 208 3145 272
rect 3049 192 3145 208
rect 3049 128 3065 192
rect 3129 128 3145 192
rect 3049 112 3145 128
rect 3049 48 3065 112
rect 3129 48 3145 112
rect 3049 32 3145 48
rect 3049 -32 3065 32
rect 3129 -32 3145 32
rect 3049 -48 3145 -32
rect 3049 -112 3065 -48
rect 3129 -112 3145 -48
rect 3049 -128 3145 -112
rect 3049 -192 3065 -128
rect 3129 -192 3145 -128
rect 3049 -208 3145 -192
rect 3049 -272 3065 -208
rect 3129 -272 3145 -208
rect 3049 -288 3145 -272
rect 3049 -352 3065 -288
rect 3129 -352 3145 -288
rect 3049 -368 3145 -352
rect 3049 -432 3065 -368
rect 3129 -432 3145 -368
rect 3049 -448 3145 -432
rect 3049 -512 3065 -448
rect 3129 -512 3145 -448
rect 3049 -528 3145 -512
rect 3049 -592 3065 -528
rect 3129 -592 3145 -528
rect 3049 -608 3145 -592
rect 3049 -672 3065 -608
rect 3129 -672 3145 -608
rect 3049 -688 3145 -672
rect 3049 -752 3065 -688
rect 3129 -752 3145 -688
rect 3049 -768 3145 -752
rect 3049 -832 3065 -768
rect 3129 -832 3145 -768
rect 3049 -848 3145 -832
rect 3049 -912 3065 -848
rect 3129 -912 3145 -848
rect 3049 -928 3145 -912
rect 3049 -992 3065 -928
rect 3129 -992 3145 -928
rect 3049 -1008 3145 -992
rect 3049 -1072 3065 -1008
rect 3129 -1072 3145 -1008
rect 3049 -1088 3145 -1072
<< properties >>
string FIXED_BBOX -3150 -1100 3050 1100
<< end >>
