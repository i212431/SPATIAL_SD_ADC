magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< nwell >>
rect 5404 4055 5574 4271
<< locali >>
rect 536 5107 10385 5124
rect 536 4569 577 5107
rect 10331 4569 10385 5107
rect 536 4549 10385 4569
rect 3906 2687 5042 4549
rect 2454 379 3931 419
rect 107 -163 3931 379
rect 2454 -3516 3931 -163
rect 2454 -3910 2511 -3516
rect 3841 -3910 3931 -3516
rect 2454 -3971 3931 -3910
<< viali >>
rect 577 4569 10331 5107
rect 2511 -3910 3841 -3516
<< metal1 >>
rect 536 5107 10385 5124
rect 536 5088 577 5107
rect 10331 5088 10385 5107
rect 536 4588 564 5088
rect 10344 4588 10385 5088
rect 536 4569 577 4588
rect 10331 4569 10385 4588
rect 536 4549 10385 4569
rect 5404 4227 5574 4271
rect 5404 4111 5431 4227
rect 5547 4111 5574 4227
rect 5404 4055 5574 4111
rect -584 2120 -144 2191
rect -584 1556 -524 2120
rect -216 1859 -144 2120
rect -216 1795 1197 1859
rect -216 1556 -144 1795
rect -584 1496 -144 1556
rect -1045 833 -144 936
rect -1045 333 -947 833
rect -255 659 -144 833
rect -255 595 620 659
rect -255 333 -144 595
rect -1045 241 -144 333
rect 2454 -3495 3931 -3433
rect 2454 -3931 2510 -3495
rect 3842 -3931 3931 -3495
rect 2454 -3971 3931 -3931
<< via1 >>
rect 564 4588 577 5088
rect 577 4588 10331 5088
rect 10331 4588 10344 5088
rect 5431 4111 5547 4227
rect -524 1556 -216 2120
rect -947 333 -255 833
rect 2510 -3516 3842 -3495
rect 2510 -3910 2511 -3516
rect 2511 -3910 3841 -3516
rect 3841 -3910 3842 -3516
rect 2510 -3931 3842 -3910
<< metal2 >>
rect -6210 11358 16896 11472
rect -6210 9142 -6119 11358
rect -4143 11322 16896 11358
rect -4143 11276 14799 11322
rect -4143 9220 -1569 11276
rect -1193 11118 14799 11276
rect -1193 9302 11876 11118
rect 13292 9302 14799 11118
rect -1193 9220 14799 9302
rect -4143 9186 14799 9220
rect 16775 9186 16896 11322
rect -4143 9142 16896 9186
rect -6210 9064 16896 9142
rect -3284 8615 13696 8753
rect -3284 8613 12073 8615
rect -3284 7037 -3177 8613
rect -1681 8365 12073 8613
rect -1681 7589 1042 8365
rect 10938 7589 12073 8365
rect -1681 7039 12073 7589
rect 13569 7039 13696 8615
rect -1681 7037 13696 7039
rect -3284 6926 13696 7037
rect 553 5124 10361 6926
rect 536 5088 10385 5124
rect 536 4588 564 5088
rect 10344 4588 10385 5088
rect 536 4549 10385 4588
rect 1009 4239 1098 4261
rect 1009 4183 1025 4239
rect 1081 4183 1098 4239
rect 1009 4161 1098 4183
rect 2589 4242 2678 4264
rect 4259 4255 5574 4271
rect 2589 4186 2605 4242
rect 2661 4186 2678 4242
rect 2589 4164 2678 4186
rect 4135 4238 5574 4255
rect 4135 4182 4147 4238
rect 4203 4182 4227 4238
rect 4283 4182 4307 4238
rect 4363 4182 4387 4238
rect 4443 4182 4467 4238
rect 4523 4182 4547 4238
rect 4603 4182 4627 4238
rect 4683 4182 4707 4238
rect 4763 4227 5574 4238
rect 4763 4182 5431 4227
rect 4135 4165 5431 4182
rect 4259 4155 5431 4165
rect 5404 4111 5431 4155
rect 5547 4111 5574 4227
rect 5404 4055 5574 4111
rect 10166 3871 13700 3950
rect 10166 3255 12039 3871
rect 13615 3255 13700 3871
rect 593 3225 674 3240
rect 593 3169 605 3225
rect 661 3169 674 3225
rect 593 3155 674 3169
rect 3591 3229 3672 3244
rect 3591 3173 3603 3229
rect 3659 3173 3672 3229
rect 10166 3206 13700 3255
rect 3591 3159 3672 3173
rect -9221 2120 -144 2191
rect -9221 1556 -524 2120
rect -216 1556 -144 2120
rect 9560 2048 11023 2119
rect -9221 1496 -144 1556
rect 1003 1633 1092 1655
rect 1003 1577 1019 1633
rect 1075 1577 1092 1633
rect 1003 1555 1092 1577
rect 2582 1632 2671 1654
rect 2582 1576 2598 1632
rect 2654 1576 2671 1632
rect 2582 1554 2671 1576
rect 9560 1432 10667 2048
rect 10963 1432 11023 2048
rect 9560 1372 11023 1432
rect 866 1289 1072 1307
rect 866 1233 901 1289
rect 957 1233 981 1289
rect 1037 1233 1072 1289
rect 866 1215 1072 1233
rect 1498 1290 1704 1308
rect 1498 1234 1533 1290
rect 1589 1234 1613 1290
rect 1669 1234 1704 1290
rect 1498 1216 1704 1234
rect -9221 833 -144 936
rect -9221 333 -947 833
rect -255 333 -144 833
rect 530 864 611 879
rect 530 808 542 864
rect 598 808 611 864
rect 530 794 611 808
rect 3531 864 3612 879
rect 3531 808 3543 864
rect 3599 808 3612 864
rect 3531 794 3612 808
rect -9221 241 -144 333
rect -9176 -401 -125 -163
rect -9176 -567 485 -401
rect -9176 -858 -125 -567
rect 864 -776 1072 -754
rect 864 -912 900 -776
rect 1036 -912 1072 -776
rect 864 -933 1072 -912
rect 1500 -775 1708 -753
rect 1500 -911 1536 -775
rect 1672 -911 1708 -775
rect 1500 -932 1708 -911
rect 2108 -1737 11865 -1636
rect 2108 -2273 10705 -1737
rect 11721 -2273 11865 -1737
rect 2108 -2389 11865 -2273
rect 2454 -3485 3931 -3433
rect 2454 -3941 2508 -3485
rect 3844 -3941 3931 -3485
rect 2454 -3971 3931 -3941
rect -3284 -5480 13696 -5334
rect -3284 -5519 12128 -5480
rect -3284 -7015 -3149 -5519
rect -1813 -6976 12128 -5519
rect 13464 -6976 13696 -5480
rect -1813 -7015 13696 -6976
rect -3284 -7161 13696 -7015
rect -6210 -7775 16896 -7596
rect -6210 -7806 2590 -7775
rect -6210 -9862 -6104 -7806
rect -4128 -9831 2590 -7806
rect 3766 -7795 16896 -7775
rect 3766 -9771 14862 -7795
rect 16678 -9771 16896 -7795
rect 3766 -9831 16896 -9771
rect -4128 -9862 16896 -9831
rect -6210 -10004 16896 -9862
<< via2 >>
rect -6119 9142 -4143 11358
rect -1569 9220 -1193 11276
rect 11876 9302 13292 11118
rect 14799 9186 16775 11322
rect -3177 7037 -1681 8613
rect 1042 7589 10938 8365
rect 12073 7039 13569 8615
rect 1025 4183 1081 4239
rect 2605 4186 2661 4242
rect 4147 4182 4203 4238
rect 4227 4182 4283 4238
rect 4307 4182 4363 4238
rect 4387 4182 4443 4238
rect 4467 4182 4523 4238
rect 4547 4182 4603 4238
rect 4627 4182 4683 4238
rect 4707 4182 4763 4238
rect 12039 3255 13615 3871
rect 605 3169 661 3225
rect 3603 3173 3659 3229
rect 1019 1577 1075 1633
rect 2598 1576 2654 1632
rect 10667 1432 10963 2048
rect 901 1233 957 1289
rect 981 1233 1037 1289
rect 1533 1234 1589 1290
rect 1613 1234 1669 1290
rect 542 808 598 864
rect 3543 808 3599 864
rect 900 -912 1036 -776
rect 1536 -911 1672 -775
rect 10705 -2273 11721 -1737
rect 2508 -3495 3844 -3485
rect 2508 -3931 2510 -3495
rect 2510 -3931 3842 -3495
rect 3842 -3931 3844 -3495
rect 2508 -3941 3844 -3931
rect -3149 -7015 -1813 -5519
rect 12128 -6976 13464 -5480
rect -6104 -9862 -4128 -7806
rect 2590 -9831 3766 -7775
rect 14862 -9771 16678 -7795
<< metal3 >>
rect -6210 11358 -4008 11474
rect -6210 9142 -6119 11358
rect -4143 9142 -4008 11358
rect -6210 9064 -4008 9142
rect -1700 11280 -1041 11472
rect -1700 9216 -1573 11280
rect -1189 9216 -1041 11280
rect -1700 9064 -1041 9216
rect 11720 11122 13486 11472
rect 11720 11118 11912 11122
rect 13256 11118 13486 11122
rect 11720 9302 11876 11118
rect 13292 9302 13486 11118
rect 11720 9298 11912 9302
rect 13256 9298 13486 9302
rect 11720 9064 13486 9298
rect 14675 11322 16896 11472
rect 14675 9186 14799 11322
rect 16775 9186 16896 11322
rect -6210 -7806 -3997 9064
rect -3284 8613 -1572 8753
rect -3284 7037 -3177 8613
rect -1681 7037 -1572 8613
rect 11984 8615 13696 8753
rect 899 8369 11049 8503
rect 899 7585 1038 8369
rect 10942 7585 11049 8369
rect 899 7473 11049 7585
rect -3284 -5519 -1572 7037
rect 11984 7039 12073 8615
rect 13569 7039 13696 8615
rect 988 4239 1120 4271
rect 988 4183 1025 4239
rect 1081 4183 1120 4239
rect 459 3225 695 3260
rect 459 3169 605 3225
rect 661 3169 695 3225
rect 459 864 695 3169
rect 988 1633 1120 4183
rect 988 1577 1019 1633
rect 1075 1577 1120 1633
rect 988 1547 1120 1577
rect 2568 4242 2700 4271
rect 2568 4186 2605 4242
rect 2661 4186 2700 4242
rect 2568 1632 2700 4186
rect 4117 4238 4797 4271
rect 4117 4182 4147 4238
rect 4203 4182 4227 4238
rect 4283 4182 4307 4238
rect 4363 4182 4387 4238
rect 4443 4182 4467 4238
rect 4523 4182 4547 4238
rect 4603 4182 4627 4238
rect 4683 4182 4707 4238
rect 4763 4182 4797 4238
rect 2568 1576 2598 1632
rect 2654 1576 2700 1632
rect 2568 1547 2700 1576
rect 3451 3229 3687 3260
rect 3451 3173 3603 3229
rect 3659 3173 3687 3229
rect 459 808 542 864
rect 598 808 695 864
rect 459 775 695 808
rect 844 1289 1094 1320
rect 844 1233 901 1289
rect 957 1233 981 1289
rect 1037 1233 1094 1289
rect 844 -776 1094 1233
rect 844 -912 900 -776
rect 1036 -912 1094 -776
rect 844 -949 1094 -912
rect 1476 1290 1726 1320
rect 1476 1234 1533 1290
rect 1589 1234 1613 1290
rect 1669 1234 1726 1290
rect 1476 -775 1726 1234
rect 3451 864 3687 3173
rect 3451 808 3543 864
rect 3599 808 3687 864
rect 3451 775 3687 808
rect 1476 -911 1536 -775
rect 1672 -911 1726 -775
rect 1476 -949 1726 -911
rect 4117 -801 4797 4182
rect 11984 3871 13696 7039
rect 11984 3255 12039 3871
rect 13615 3255 13696 3871
rect 10624 2052 11023 2119
rect 10624 2048 10703 2052
rect 10927 2048 11023 2052
rect 10624 1432 10667 2048
rect 10963 1432 11023 2048
rect 10624 1428 10703 1432
rect 10927 1428 11023 1432
rect 10624 1372 11023 1428
rect 4117 -2945 4180 -801
rect 4724 -2945 4797 -801
rect 10524 -1733 11865 -1636
rect 10524 -1737 10741 -1733
rect 11685 -1737 11865 -1733
rect 10524 -2273 10705 -1737
rect 11721 -2273 11865 -1737
rect 10524 -2277 10741 -2273
rect 11685 -2277 11865 -2273
rect 10524 -2389 11865 -2277
rect 4117 -3017 4797 -2945
rect -3284 -7015 -3149 -5519
rect -1813 -7015 -1572 -5519
rect -3284 -7161 -1572 -7015
rect 2454 -3485 3931 -3433
rect 2454 -3941 2508 -3485
rect 3844 -3941 3931 -3485
rect -6210 -9862 -6104 -7806
rect -4128 -9862 -3997 -7806
rect -6210 -10004 -3997 -9862
rect 2454 -7775 3931 -3941
rect 11984 -5480 13696 3255
rect 11984 -6976 12128 -5480
rect 13464 -6976 13696 -5480
rect 11984 -7161 13696 -6976
rect 2454 -9831 2590 -7775
rect 3766 -9831 3931 -7775
rect 2454 -10004 3931 -9831
rect 14675 -7795 16896 9186
rect 14675 -9771 14862 -7795
rect 16678 -9771 16896 -7795
rect 14675 -10004 16896 -9771
<< via3 >>
rect -1573 11276 -1189 11280
rect -1573 9220 -1569 11276
rect -1569 9220 -1193 11276
rect -1193 9220 -1189 11276
rect -1573 9216 -1189 9220
rect 11912 11118 13256 11122
rect 11912 9302 13256 11118
rect 11912 9298 13256 9302
rect 1038 8365 10942 8369
rect 1038 7589 1042 8365
rect 1042 7589 10938 8365
rect 10938 7589 10942 8365
rect 1038 7585 10942 7589
rect 10703 2048 10927 2052
rect 10703 1432 10927 2048
rect 10703 1428 10927 1432
rect 4180 -2945 4724 -801
rect 10741 -1737 11685 -1733
rect 10741 -2273 11685 -1737
rect 10741 -2277 11685 -2273
<< metal4 >>
rect -1700 11280 -1041 11472
rect -1700 9216 -1573 11280
rect -1189 9216 -1041 11280
rect -1700 5103 -1041 9216
rect 11720 11122 13486 11472
rect 11720 9298 11912 11122
rect 13256 9298 13486 11122
rect 899 8369 11049 8503
rect 899 7585 1038 8369
rect 10942 7585 11049 8369
rect 899 6726 11049 7585
rect 899 5452 11084 6726
rect 11720 5102 13486 9298
rect 10624 2052 12031 2121
rect 10624 1428 10703 2052
rect 10927 1428 12031 2052
rect 10624 995 12031 1428
rect 10624 61 21004 995
rect 4117 -801 8769 -674
rect 4117 -2945 4180 -801
rect 4724 -2945 8769 -801
rect 4117 -3017 8769 -2945
rect 10524 -920 21004 61
rect 10524 -1636 11023 -920
rect 11612 -1424 21004 -920
rect 10524 -1733 11865 -1636
rect 10524 -2277 10741 -1733
rect 11685 -2277 11865 -1733
rect 10524 -2389 11865 -2277
rect 10524 -4915 11023 -2389
use CurrentMirror_layout  CurrentMirror_layout_0
timestamp 1667803582
transform 1 0 634 0 1 -2505
box -553 -441 2226 2534
use DiffPair_layout  DiffPair_layout_0
timestamp 1667803582
transform 1 0 462 0 1 701
box -415 -553 3823 1603
use PMOS2  PMOS2_0
timestamp 1667803582
transform 1 0 4139 0 1 1699
box 509 -1491 6581 3083
use PMOS_Load  PMOS_Load_0
timestamp 1667803582
transform 1 0 490 0 1 3052
box -508 -541 3903 1749
use sky130_fd_pr__cap_mim_m3_1_N3PKNJ  sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0
timestamp 1667803582
transform 1 0 8671 0 1 6190
box -3150 -1100 3149 1100
use sky130_fd_pr__cap_mim_m3_1_N3PKNJ  sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1
timestamp 1667803582
transform -1 0 2036 0 1 6190
box -3150 -1100 3149 1100
use sky130_fd_pr__cap_mim_m3_1_TQVBRR  sky130_fd_pr__cap_mim_m3_1_TQVBRR_0
timestamp 1667803582
transform 1 0 8075 0 1 -2427
box -2550 -2500 2549 2500
<< labels >>
flabel metal2 s -8791 531 -8791 531 0 FreeSans 3125 0 0 0 VN
port 1 nsew
flabel metal2 s -8568 1903 -8568 1903 0 FreeSans 3125 0 0 0 VP
port 2 nsew
flabel metal2 s -8852 -591 -8852 -591 0 FreeSans 3125 0 0 0 IBIAS
port 3 nsew
flabel metal3 s 5485 7900 5485 7900 0 FreeSans 9375 0 0 0 VDD
port 4 nsew
flabel metal2 s 5268 10390 5268 10390 0 FreeSans 9375 0 0 0 VSS
port 5 nsew
flabel metal4 s 19494 -84 19494 -84 0 FreeSans 9375 0 0 0 VO
port 6 nsew
<< end >>
