* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130B

.subckt sky130_fd_sc_hd__clkbuf_4 X A VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=9.1e+11p pd=7.82e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=3.801e+11p pd=4.33e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_LZABJ9 a_n73_n64# a_n33_n161# li_n175_n248# a_15_n64#
+ w_n211_n284#
X0 a_15_n64# a_n33_n161# a_n73_n64# w_n211_n284# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_LTABJ9 a_n33_n461# a_15_n364# li_n175_n548# w_n211_n584#
+ a_n73_n364#
X0 a_15_n364# a_n33_n461# a_n73_n364# w_n211_n584# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_RB5HKB a_15_n131# a_n175_n243# a_n33_91# li_n175_n243#
+ a_n73_n131#
X0 a_15_n131# a_n33_91# a_n73_n131# a_n175_n243# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_6H5H3D li_n175_n343# a_n33_191# a_n73_n231# a_15_n231#
+ a_n175_n343#
X0 a_15_n231# a_n33_191# a_n73_n231# a_n175_n343# sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_LDKBCP a_n73_n81# a_n175_n193# li_n175_n193# a_n33_41#
+ a_15_n81#
X0 a_15_n81# a_n33_41# a_n73_n81# a_n175_n193# sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
.ends

.subckt COMPA VOUTP VDD VOUTN VINN CLK VINP VSS
Xsky130_fd_pr__pfet_01v8_LZABJ9_3 VDD CLK sky130_fd_pr__pfet_01v8_LZABJ9_5/li_n175_n248#
+ m1_113_808# VDD sky130_fd_pr__pfet_01v8_LZABJ9
Xsky130_fd_pr__pfet_01v8_LZABJ9_5 m1_113_808# m1_757_1008# sky130_fd_pr__pfet_01v8_LZABJ9_5/li_n175_n248#
+ VDD VDD sky130_fd_pr__pfet_01v8_LZABJ9
Xsky130_fd_pr__pfet_01v8_LZABJ9_4 m1_541_888# CLK sky130_fd_pr__pfet_01v8_LZABJ9_5/li_n175_n248#
+ VDD VDD sky130_fd_pr__pfet_01v8_LZABJ9
Xsky130_fd_pr__pfet_01v8_LTABJ9_0 m1_757_1008# VOUTN sky130_fd_pr__pfet_01v8_LZABJ9_2/li_n175_n248#
+ VDD VDD sky130_fd_pr__pfet_01v8_LTABJ9
Xsky130_fd_pr__pfet_01v8_LTABJ9_1 m1_113_808# VDD sky130_fd_pr__pfet_01v8_LZABJ9_5/li_n175_n248#
+ VDD VOUTP sky130_fd_pr__pfet_01v8_LTABJ9
Xsky130_fd_pr__nfet_01v8_RB5HKB_0 m1_383_104# VSS CLK sky130_fd_pr__nfet_01v8_RB5HKB_0/li_n175_n243#
+ VSS sky130_fd_pr__nfet_01v8_RB5HKB
Xsky130_fd_pr__nfet_01v8_6H5H3D_0 sky130_fd_pr__nfet_01v8_6H5H3D_1/li_n175_n343# m1_757_1008#
+ VSS VOUTN VSS sky130_fd_pr__nfet_01v8_6H5H3D
Xsky130_fd_pr__pfet_01v8_LZABJ9_0 VDD CLK sky130_fd_pr__pfet_01v8_LZABJ9_2/li_n175_n248#
+ m1_1362_377# VDD sky130_fd_pr__pfet_01v8_LZABJ9
Xsky130_fd_pr__nfet_01v8_6H5H3D_1 sky130_fd_pr__nfet_01v8_6H5H3D_1/li_n175_n343# VINN
+ m1_1362_377# m1_383_104# VSS sky130_fd_pr__nfet_01v8_6H5H3D
Xsky130_fd_pr__nfet_01v8_LDKBCP_0 m1_757_1008# VSS sky130_fd_pr__nfet_01v8_RB5HKB_0/li_n175_n243#
+ m1_113_808# m1_1362_377# sky130_fd_pr__nfet_01v8_LDKBCP
Xsky130_fd_pr__pfet_01v8_LZABJ9_1 m1_757_1008# CLK sky130_fd_pr__pfet_01v8_LZABJ9_2/li_n175_n248#
+ VDD VDD sky130_fd_pr__pfet_01v8_LZABJ9
Xsky130_fd_pr__nfet_01v8_LDKBCP_1 m1_541_888# VSS sky130_fd_pr__nfet_01v8_RB5HKB_0/li_n175_n243#
+ m1_757_1008# m1_113_808# sky130_fd_pr__nfet_01v8_LDKBCP
Xsky130_fd_pr__nfet_01v8_6H5H3D_2 sky130_fd_pr__nfet_01v8_6H5H3D_3/li_n175_n343# VINP
+ m1_383_104# m1_541_888# VSS sky130_fd_pr__nfet_01v8_6H5H3D
Xsky130_fd_pr__pfet_01v8_LZABJ9_2 VDD m1_113_808# sky130_fd_pr__pfet_01v8_LZABJ9_2/li_n175_n248#
+ m1_757_1008# VDD sky130_fd_pr__pfet_01v8_LZABJ9
Xsky130_fd_pr__nfet_01v8_6H5H3D_3 sky130_fd_pr__nfet_01v8_6H5H3D_3/li_n175_n343# m1_113_808#
+ VOUTP VSS VSS sky130_fd_pr__nfet_01v8_6H5H3D
.ends

.subckt sky130_fd_sc_hd__clkinv_16 Y A VGND VPWR VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.0605e+12p pd=1.261e+07u as=1.0059e+12p ps=1.151e+07u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.515e+12p pd=3.103e+07u as=3.655e+12p ps=3.331e+07u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_52DJHB a_n129_n500# a_63_n500# a_15_n597# a_n81_531#
+ a_n177_n597# w_n257_n600# a_n33_n500# a_159_n500# a_111_531# a_n221_n500#
X0 a_n33_n500# a_n81_531# a_n129_n500# w_n257_n600# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X1 a_159_n500# a_111_531# a_63_n500# w_n257_n600# sky130_fd_pr__pfet_01v8 ad=1.55e+12p pd=1.062e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X2 a_63_n500# a_15_n597# a_n33_n500# w_n257_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3 a_n129_n500# a_n177_n597# a_n221_n500# w_n257_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.55e+12p ps=1.062e+07u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_JRYMCH a_n33_n250# a_n81_272# a_159_n250# a_15_n338#
+ a_n177_n338# a_n221_n250# a_n129_n250# a_63_n250# a_111_272# VSUBS
X0 a_n129_n250# a_n177_n338# a_n221_n250# VSUBS sky130_fd_pr__nfet_01v8 ad=8.25e+11p pd=5.66e+06u as=7.75e+11p ps=5.62e+06u w=2.5e+06u l=150000u
X1 a_n33_n250# a_n81_272# a_n129_n250# VSUBS sky130_fd_pr__nfet_01v8 ad=8.25e+11p pd=5.66e+06u as=0p ps=0u w=2.5e+06u l=150000u
X2 a_159_n250# a_111_272# a_63_n250# VSUBS sky130_fd_pr__nfet_01v8 ad=7.75e+11p pd=5.62e+06u as=8.25e+11p ps=5.66e+06u w=2.5e+06u l=150000u
X3 a_63_n250# a_15_n338# a_n33_n250# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
.ends

.subckt T_Gate B A CLKB VDD sky130_fd_sc_hd__clkinv_16_0/A VSS
Xsky130_fd_sc_hd__clkinv_16_0 CLKB sky130_fd_sc_hd__clkinv_16_0/A VSS VDD VSS VDD
+ sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__pfet_01v8_52DJHB_0 A A CLKB CLKB CLKB VDD B B CLKB B sky130_fd_pr__pfet_01v8_52DJHB
Xsky130_fd_pr__nfet_01v8_JRYMCH_0 B sky130_fd_sc_hd__clkinv_16_0/A B sky130_fd_sc_hd__clkinv_16_0/A
+ sky130_fd_sc_hd__clkinv_16_0/A B A A sky130_fd_sc_hd__clkinv_16_0/A VSS sky130_fd_pr__nfet_01v8_JRYMCH
.ends

.subckt sky130_fd_pr__nfet_01v8_H73VBR a_n33_n250# a_n81_272# a_159_n250# a_15_n338#
+ a_n177_n338# a_n221_n250# a_n129_n250# a_63_n250# a_n323_n424# a_111_272#
X0 a_n129_n250# a_n177_n338# a_n221_n250# a_n323_n424# sky130_fd_pr__nfet_01v8 ad=8.25e+11p pd=5.66e+06u as=7.75e+11p ps=5.62e+06u w=2.5e+06u l=150000u
X1 a_n33_n250# a_n81_272# a_n129_n250# a_n323_n424# sky130_fd_pr__nfet_01v8 ad=8.25e+11p pd=5.66e+06u as=0p ps=0u w=2.5e+06u l=150000u
X2 a_159_n250# a_111_272# a_63_n250# a_n323_n424# sky130_fd_pr__nfet_01v8 ad=7.75e+11p pd=5.62e+06u as=8.25e+11p ps=5.66e+06u w=2.5e+06u l=150000u
X3 a_63_n250# a_15_n338# a_n33_n250# a_n323_n424# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MJDHVK m3_n2950_n2900# c1_n2850_n2800#
X0 c1_n2850_n2800# m3_n2950_n2900# sky130_fd_pr__cap_mim_m3_1 l=2.8e+07u w=2.8e+07u
.ends

.subckt Subtractor_Mag VGND PH2 VOUT T_Gate_1/sky130_fd_sc_hd__clkinv_16_0/A T_Gate_0/B
+ T_Gate_0/A T_Gate_1/VDD T_Gate_1/B VSUBS
XT_Gate_0 T_Gate_0/B T_Gate_0/A T_Gate_0/CLKB T_Gate_1/VDD T_Gate_1/sky130_fd_sc_hd__clkinv_16_0/A
+ VSUBS T_Gate
XT_Gate_1 T_Gate_1/B VOUT T_Gate_1/CLKB T_Gate_1/VDD T_Gate_1/sky130_fd_sc_hd__clkinv_16_0/A
+ VSUBS T_Gate
Xsky130_fd_pr__nfet_01v8_H73VBR_0 T_Gate_0/B PH2 T_Gate_0/B PH2 PH2 T_Gate_0/B VGND
+ VGND VSUBS PH2 sky130_fd_pr__nfet_01v8_H73VBR
Xsky130_fd_pr__cap_mim_m3_1_MJDHVK_0 T_Gate_0/B VOUT sky130_fd_pr__cap_mim_m3_1_MJDHVK
.ends

.subckt sky130_fd_pr__nfet_01v8_RC9KLY a_50_n1050# a_n50_n1076# a_n108_n1050# VSUBS
X0 a_50_n1050# a_n50_n1076# a_n108_n1050# VSUBS sky130_fd_pr__nfet_01v8 ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=500000u
.ends

.subckt CurrentMirror_layout D3 S D1 D2
Xsky130_fd_pr__nfet_01v8_RC9KLY_1 D3 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_2 S D1 D3 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_3 S D1 D1 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_4 S D1 D3 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_5 D1 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_6 S D1 D2 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_7 D3 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_8 S D1 D3 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_9 D2 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_0 D3 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
.ends

.subckt sky130_fd_pr__nfet_01v8_6YBK2C a_50_n500# a_n50_n526# a_n108_n500# VSUBS
X0 a_50_n500# a_n50_n526# a_n108_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt DiffPair_layout G1 G2 D2 S D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
Xsky130_fd_pr__nfet_01v8_6YBK2C_10 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_11 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_12 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_13 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_14 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_15 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_16 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_17 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_18 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_19 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_0 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_1 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_2 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_3 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_4 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_5 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_6 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_7 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_8 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_9 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_EEU9S7 w_n144_n662# a_50_n600# a_n50_n626# a_n108_n600#
X0 a_50_n600# a_n50_n626# a_n108_n600# w_n144_n662# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
.ends

.subckt PMOS_Load D2 D1 S
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_0 S D1 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_1 S S D1 D2 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_2 S D2 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_10 S S D1 D1 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_3 S S D1 D1 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_11 S D2 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_4 S D1 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_12 S S D1 D2 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_5 S S D1 D2 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_13 S D1 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_6 S D2 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_7 S S D1 D1 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_14 S S D1 D1 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_8 S D1 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_15 S D2 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_9 S S D1 D2 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_16 S S D1 D2 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_17 S D1 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_18 S S D1 D1 sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_19 S D2 D1 S sky130_fd_pr__pfet_01v8_lvt_EEU9S7
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_TQVBRR m3_n2550_n2500# c1_n2450_n2400#
X0 c1_n2450_n2400# m3_n2550_n2500# sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.4e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_N3PKNJ c1_n3050_n1000# m3_n3150_n1100#
X0 c1_n3050_n1000# m3_n3150_n1100# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_WFBLZ7 a_50_n1420# a_n50_n1446# w_n144_n1482#
+ a_n108_n1420#
X0 a_50_n1420# a_n50_n1446# a_n108_n1420# w_n144_n1482# sky130_fd_pr__pfet_01v8_lvt ad=4.118e+12p pd=2.898e+07u as=4.118e+12p ps=2.898e+07u w=1.42e+07u l=500000u
.ends

.subckt PMOS2 S D G
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_19 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_0 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_1 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_2 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_3 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_4 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_5 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_6 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_7 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_8 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_9 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_20 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_10 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_21 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_11 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_22 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_12 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_23 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_13 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_24 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_14 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_15 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_16 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_17 D G S S sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_18 S G S D sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
.ends

.subckt OpampM VN VP IBIAS VDD VSS VO
XCurrentMirror_layout_0 VO VSS IBIAS DiffPair_layout_0/S CurrentMirror_layout
XDiffPair_layout_0 VN VP PMOS2_0/G DiffPair_layout_0/S PMOS_Load_0/D1 VSS DiffPair_layout
XPMOS_Load_0 PMOS2_0/G PMOS_Load_0/D1 VDD PMOS_Load
Xsky130_fd_pr__cap_mim_m3_1_TQVBRR_0 VO PMOS2_0/G sky130_fd_pr__cap_mim_m3_1_TQVBRR
Xsky130_fd_pr__cap_mim_m3_1_N3PKNJ_0 VDD VSS sky130_fd_pr__cap_mim_m3_1_N3PKNJ
Xsky130_fd_pr__cap_mim_m3_1_N3PKNJ_1 VDD VSS sky130_fd_pr__cap_mim_m3_1_N3PKNJ
XPMOS2_0 VDD VO PMOS2_0/G PMOS2
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_4RKXMF m3_n2950_n2900# c1_n2850_n2800#
X0 c1_n2850_n2800# m3_n2950_n2900# sky130_fd_pr__cap_mim_m3_1 l=2.8e+07u w=2.8e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_FR7DL7 a_n33_n250# a_n81_272# a_159_n250# a_15_n338#
+ a_n177_n338# a_n221_n250# a_n129_n250# a_63_n250# a_n323_n424# a_111_272#
X0 a_n129_n250# a_n177_n338# a_n221_n250# a_n323_n424# sky130_fd_pr__nfet_01v8 ad=8.25e+11p pd=5.66e+06u as=7.75e+11p ps=5.62e+06u w=2.5e+06u l=150000u
X1 a_n33_n250# a_n81_272# a_n129_n250# a_n323_n424# sky130_fd_pr__nfet_01v8 ad=8.25e+11p pd=5.66e+06u as=0p ps=0u w=2.5e+06u l=150000u
X2 a_159_n250# a_111_272# a_63_n250# a_n323_n424# sky130_fd_pr__nfet_01v8 ad=7.75e+11p pd=5.62e+06u as=8.25e+11p ps=5.66e+06u w=2.5e+06u l=150000u
X3 a_63_n250# a_15_n338# a_n33_n250# a_n323_n424# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
.ends

.subckt co VDD VREF VIN VOUT PH1 PH2 VSS
XT_Gate_0 T_Gate_0/B VIN T_Gate_0/CLKB VDD PH1 VSS T_Gate
XT_Gate_1 VOUT T_Gate_1/A T_Gate_1/CLKB VDD PH2 VSS T_Gate
Xsky130_fd_pr__cap_mim_m3_1_4RKXMF_0 T_Gate_1/A T_Gate_0/B sky130_fd_pr__cap_mim_m3_1_4RKXMF
Xsky130_fd_pr__nfet_01v8_FR7DL7_0 VREF PH1 VREF PH1 PH1 VREF T_Gate_1/A T_Gate_1/A
+ VSS PH1 sky130_fd_pr__nfet_01v8_FR7DL7
Xsky130_fd_pr__nfet_01v8_FR7DL7_1 VREF PH2 VREF PH2 PH2 VREF T_Gate_0/B T_Gate_0/B
+ VSS PH2 sky130_fd_pr__nfet_01v8_FR7DL7
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_D7CHNQ c1_n1550_n1500# m3_n1650_n1600#
X0 c1_n1550_n1500# m3_n1650_n1600# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
.ends

.subckt Integrator_n co_0/VIN co_0/PH1 co_0/VREF co_0/PH2 OpampM_0/IBIAS co_0/VDD
+ VSUBS OpampM_0/VO
XOpampM_0 co_0/VOUT co_0/VREF OpampM_0/IBIAS co_0/VDD VSUBS OpampM_0/VO OpampM
Xco_0 co_0/VDD co_0/VREF co_0/VIN co_0/VOUT co_0/PH1 co_0/PH2 VSUBS co
Xsky130_fd_pr__cap_mim_m3_1_D7CHNQ_0 co_0/VOUT OpampM_0/VO sky130_fd_pr__cap_mim_m3_1_D7CHNQ
.ends

.subckt sky130_fd_sc_hd__bufbuf_16 A X VGND VPWR VNB VPB
X0 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.16e+12p pd=2.032e+07u as=3.76e+12p ps=3.552e+07u w=1e+06u l=150000u
X1 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.404e+12p pd=1.472e+07u as=2.444e+12p ps=2.572e+07u w=650000u l=150000u
X2 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X3 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X4 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X7 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X36 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X45 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X47 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X51 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A X VGND VPWR VNB VPB
X0 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=6.517e+11p ps=5.37e+06u w=820000u l=500000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=4.027e+11p pd=3.97e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X7 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt Delay_Block VOUT VIN VSS VDD
Xsky130_fd_sc_hd__clkdlybuf4s50_1_0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/X VOUT VSS
+ VDD VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_1 VIN sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS VDD
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_2 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
.ends

.subckt sky130_fd_pr__nfet_01v8_WWN8PW a_n33_n250# a_n81_272# a_159_n250# a_15_n338#
+ a_n177_n338# a_n221_n250# a_n129_n250# a_63_n250# a_111_272# VSUBS
X0 a_n129_n250# a_n177_n338# a_n221_n250# VSUBS sky130_fd_pr__nfet_01v8 ad=8.25e+11p pd=5.66e+06u as=7.75e+11p ps=5.62e+06u w=2.5e+06u l=150000u
X1 a_n33_n250# a_n81_272# a_n129_n250# VSUBS sky130_fd_pr__nfet_01v8 ad=8.25e+11p pd=5.66e+06u as=0p ps=0u w=2.5e+06u l=150000u
X2 a_159_n250# a_111_272# a_63_n250# VSUBS sky130_fd_pr__nfet_01v8 ad=7.75e+11p pd=5.62e+06u as=8.25e+11p ps=5.66e+06u w=2.5e+06u l=150000u
X3 a_63_n250# a_15_n338# a_n33_n250# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
.ends

.subckt DAC VREF_P VREF_N VOUT VIN VDD VSS
Xsky130_fd_sc_hd__clkinv_16_0 sky130_fd_sc_hd__clkinv_16_0/Y VIN VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__pfet_01v8_52DJHB_0 VREF_N VREF_N sky130_fd_sc_hd__clkinv_16_0/Y sky130_fd_sc_hd__clkinv_16_0/Y
+ sky130_fd_sc_hd__clkinv_16_0/Y VDD VOUT VOUT sky130_fd_sc_hd__clkinv_16_0/Y VOUT
+ sky130_fd_pr__pfet_01v8_52DJHB
Xsky130_fd_pr__pfet_01v8_52DJHB_1 VREF_P VREF_P VIN VIN VIN VDD VOUT VOUT VIN VOUT
+ sky130_fd_pr__pfet_01v8_52DJHB
Xsky130_fd_pr__nfet_01v8_WWN8PW_0 VOUT sky130_fd_sc_hd__clkinv_16_0/Y VOUT sky130_fd_sc_hd__clkinv_16_0/Y
+ sky130_fd_sc_hd__clkinv_16_0/Y VOUT VREF_P VREF_P sky130_fd_sc_hd__clkinv_16_0/Y
+ VSS sky130_fd_pr__nfet_01v8_WWN8PW
Xsky130_fd_pr__nfet_01v8_WWN8PW_1 VOUT VIN VOUT VIN VIN VOUT VREF_N VREF_N VIN VSS
+ sky130_fd_pr__nfet_01v8_WWN8PW
.ends

.subckt sky130_fd_sc_hd__nor2_1 B Y A VGND VPWR VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 Y A VGND VPWR VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=4.536e+11p ps=4.44e+06u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.197e+11p pd=1.41e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt NOCFINAL PH1 CLK VDD PH2 sky130_fd_sc_hd__clkdlybuf4s50_1_0/X VSS
Xsky130_fd_sc_hd__clkdlybuf4s50_1_0 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_0/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_1 sky130_fd_sc_hd__nor2_1_1/Y PH2 VSS VDD VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nor2_1_0 PH2 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__nor2_1_0/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 PH1 sky130_fd_sc_hd__nor2_1_1/Y CLK VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__nor2_1_0/A CLK VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPWR VGND VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=7.492e+11p ps=8.11e+06u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.02105e+12p pd=9.61e+06u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt TOP2nn VDD SD_IN_1 SD_DOUT_1 VQ Integrator_n_0/OpampM_0/IBIAS Subtractor_Mag_0/VOUT
+ CLK COMPA_0/VINN VSS
XCOMPA_0 COMPA_0/VOUTP VDD COMPA_0/VOUTN COMPA_0/VINN CLK COMPA_0/VINP VSS COMPA
XSubtractor_Mag_0 COMPA_0/VINN Subtractor_Mag_1/PH2 Subtractor_Mag_0/VOUT sky130_fd_sc_hd__bufbuf_16_1/X
+ Subtractor_Mag_0/T_Gate_0/B COMPA_0/VINP VDD DAC_0/VOUT VSS Subtractor_Mag
XSubtractor_Mag_1 VQ Subtractor_Mag_1/PH2 Subtractor_Mag_1/VOUT sky130_fd_sc_hd__bufbuf_16_1/X
+ Subtractor_Mag_1/T_Gate_0/B DAC_0/VOUT VDD SD_IN_1 VSS Subtractor_Mag
XIntegrator_n_0 Subtractor_Mag_1/VOUT Subtractor_Mag_1/PH2 COMPA_0/VINN sky130_fd_sc_hd__bufbuf_16_1/X
+ Integrator_n_0/OpampM_0/IBIAS VDD VSS COMPA_0/VINP Integrator_n
Xsky130_fd_sc_hd__bufbuf_16_0 sky130_fd_sc_hd__dfxtp_1_0/Q SD_DOUT_1 VSS VDD VSS VDD
+ sky130_fd_sc_hd__bufbuf_16
XDelay_Block_0 Delay_Block_0/VOUT CLK VSS VDD Delay_Block
Xsky130_fd_sc_hd__bufbuf_16_1 NOCFINAL_0/PH2 sky130_fd_sc_hd__bufbuf_16_1/X VSS VDD
+ VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_2 NOCFINAL_0/PH1 Subtractor_Mag_1/PH2 VSS VDD VSS VDD
+ sky130_fd_sc_hd__bufbuf_16
XDAC_0 VDD VSS DAC_0/VOUT SD_DOUT_1 VDD VSS DAC
XNOCFINAL_0 NOCFINAL_0/PH1 CLK VDD NOCFINAL_0/PH2 NOCFINAL_0/PH1 VSS NOCFINAL
Xsky130_fd_sc_hd__dfxtp_1_0 sky130_fd_sc_hd__dfxtp_1_0/Q Delay_Block_0/VOUT COMPA_0/VOUTP
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
.ends

.subckt TOP1nn SD_IN_1 SD_DOUT_1 Integrator_n_0/OpampM_0/IBIAS Subtractor_Mag_0/VOUT
+ CLK COMPA_0/VINN VSS VDD
XCOMPA_0 COMPA_0/VOUTP VDD COMPA_0/VOUTN COMPA_0/VINN CLK COMPA_0/VINP VSS COMPA
XSubtractor_Mag_0 COMPA_0/VINN Subtractor_Mag_1/PH2 Subtractor_Mag_0/VOUT sky130_fd_sc_hd__bufbuf_16_1/X
+ Subtractor_Mag_0/T_Gate_0/B COMPA_0/VINP VDD DAC_0/VOUT VSS Subtractor_Mag
XSubtractor_Mag_1 COMPA_0/VINN Subtractor_Mag_1/PH2 Subtractor_Mag_1/VOUT sky130_fd_sc_hd__bufbuf_16_1/X
+ Subtractor_Mag_1/T_Gate_0/B DAC_0/VOUT VDD SD_IN_1 VSS Subtractor_Mag
XIntegrator_n_0 Subtractor_Mag_1/VOUT Subtractor_Mag_1/PH2 COMPA_0/VINN sky130_fd_sc_hd__bufbuf_16_1/X
+ Integrator_n_0/OpampM_0/IBIAS VDD VSS COMPA_0/VINP Integrator_n
Xsky130_fd_sc_hd__bufbuf_16_0 sky130_fd_sc_hd__dfxtp_1_0/Q SD_DOUT_1 VSS VDD VSS VDD
+ sky130_fd_sc_hd__bufbuf_16
XDelay_Block_0 Delay_Block_0/VOUT CLK VSS VDD Delay_Block
Xsky130_fd_sc_hd__bufbuf_16_1 NOCFINAL_0/PH2 sky130_fd_sc_hd__bufbuf_16_1/X VSS VDD
+ VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_2 NOCFINAL_0/PH1 Subtractor_Mag_1/PH2 VSS VDD VSS VDD
+ sky130_fd_sc_hd__bufbuf_16
XDAC_0 VDD VSS DAC_0/VOUT SD_DOUT_1 VDD VSS DAC
XNOCFINAL_0 NOCFINAL_0/PH1 CLK VDD NOCFINAL_0/PH2 NOCFINAL_0/PH1 VSS NOCFINAL
Xsky130_fd_sc_hd__dfxtp_1_0 sky130_fd_sc_hd__dfxtp_1_0/Q Delay_Block_0/VOUT COMPA_0/VOUTP
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
.ends

.subckt TOP1234 IBIAS VDD VREF SD_IN_1 SD_DOUT_1 SD_DOUT_2 SD_IN_2 SD_IN_3 SD_DOUT_3
+ SD_IN_4 SD_DOUT_4 CLK VSS
Xsky130_fd_sc_hd__clkbuf_4_0 TOP2nn_2/CLK CLK VDD VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XTOP2nn_0 VDD SD_IN_2 SD_DOUT_2 TOP2nn_0/VQ IBIAS TOP2nn_1/VQ TOP2nn_2/CLK VREF VSS
+ TOP2nn
XTOP2nn_1 VDD SD_IN_3 TOP2nn_1/SD_DOUT_1 TOP2nn_1/VQ IBIAS TOP2nn_2/VQ TOP2nn_2/CLK
+ VREF VSS TOP2nn
XTOP2nn_2 VDD SD_IN_4 SD_DOUT_4 TOP2nn_2/VQ IBIAS TOP2nn_2/Subtractor_Mag_0/VOUT TOP2nn_2/CLK
+ VREF VSS TOP2nn
XTOP1nn_0 SD_IN_1 SD_DOUT_1 IBIAS TOP2nn_0/VQ TOP2nn_2/CLK VREF VSS VDD TOP1nn
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XTOP1234_0 TOP1234_0/IBIAS TOP1234_0/VDD TOP1234_0/VREF TOP1234_0/SD_IN_1 TOP1234_0/SD_DOUT_1
+ TOP1234_0/SD_DOUT_2 TOP1234_0/SD_IN_2 TOP1234_0/SD_IN_3 TOP1234_0/SD_DOUT_3 TOP1234_0/SD_IN_4
+ TOP1234_0/SD_DOUT_4 TOP1234_0/CLK VSUBS TOP1234
XCOMPA_0 COMPA_0/VOUTP COMPA_0/VDD COMPA_0/VOUTN COMPA_0/VINN COMPA_0/CLK COMPA_0/VINP
+ VSUBS COMPA
.ends

