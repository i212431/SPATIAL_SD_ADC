magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< pwell >>
rect -553 2308 2226 2534
rect -553 -217 -260 2308
rect 1933 -217 2226 2308
rect -553 -439 2226 -217
rect -553 -441 -260 -439
<< psubdiff >>
rect -527 2470 2200 2508
rect -527 2368 98 2470
rect 1832 2368 2200 2470
rect -527 2334 2200 2368
rect -527 2117 -286 2334
rect -289 111 -286 2117
rect -527 -243 -286 111
rect 1959 1980 2200 2334
rect 2197 -26 2200 1980
rect 1959 -243 2200 -26
rect -527 -277 2200 -243
rect -527 -379 41 -277
rect 1775 -379 2200 -277
rect -527 -413 2200 -379
rect -527 -415 -286 -413
<< psubdiffcont >>
rect 98 2368 1832 2470
rect -527 111 -289 2117
rect 1959 -26 2197 1980
rect 41 -379 1775 -277
<< poly >>
rect 58 2244 1580 2258
rect 58 2210 84 2244
rect 118 2210 152 2244
rect 186 2210 220 2244
rect 254 2210 288 2244
rect 322 2210 356 2244
rect 390 2210 424 2244
rect 458 2210 492 2244
rect 526 2210 560 2244
rect 594 2210 628 2244
rect 662 2210 696 2244
rect 730 2210 764 2244
rect 798 2210 832 2244
rect 866 2210 900 2244
rect 934 2210 968 2244
rect 1002 2210 1036 2244
rect 1070 2210 1104 2244
rect 1138 2210 1172 2244
rect 1206 2210 1240 2244
rect 1274 2210 1308 2244
rect 1342 2210 1376 2244
rect 1410 2210 1444 2244
rect 1478 2210 1512 2244
rect 1546 2210 1580 2244
rect 58 2194 1580 2210
rect 58 2152 158 2194
rect 216 2152 316 2194
rect 374 2152 474 2194
rect 532 2152 632 2194
rect 690 2152 790 2194
rect 848 2152 948 2194
rect 1006 2152 1106 2194
rect 1164 2152 1264 2194
rect 1322 2152 1422 2194
rect 1480 2152 1580 2194
rect 58 -42 158 0
rect 216 -42 316 0
rect 374 -42 474 0
rect 532 -42 632 0
rect 690 -42 790 0
rect 848 -42 948 0
rect 1006 -42 1106 0
rect 1164 -42 1264 0
rect 1322 -42 1422 0
rect 1480 -42 1580 0
rect 58 -56 1580 -42
rect 58 -90 84 -56
rect 118 -90 152 -56
rect 186 -90 220 -56
rect 254 -90 288 -56
rect 322 -90 356 -56
rect 390 -90 424 -56
rect 458 -90 492 -56
rect 526 -90 560 -56
rect 594 -90 628 -56
rect 662 -90 696 -56
rect 730 -90 764 -56
rect 798 -90 832 -56
rect 866 -90 900 -56
rect 934 -90 968 -56
rect 1002 -90 1036 -56
rect 1070 -90 1104 -56
rect 1138 -90 1172 -56
rect 1206 -90 1240 -56
rect 1274 -90 1308 -56
rect 1342 -90 1376 -56
rect 1410 -90 1444 -56
rect 1478 -90 1512 -56
rect 1546 -90 1580 -56
rect 58 -106 1580 -90
<< polycont >>
rect 84 2210 118 2244
rect 152 2210 186 2244
rect 220 2210 254 2244
rect 288 2210 322 2244
rect 356 2210 390 2244
rect 424 2210 458 2244
rect 492 2210 526 2244
rect 560 2210 594 2244
rect 628 2210 662 2244
rect 696 2210 730 2244
rect 764 2210 798 2244
rect 832 2210 866 2244
rect 900 2210 934 2244
rect 968 2210 1002 2244
rect 1036 2210 1070 2244
rect 1104 2210 1138 2244
rect 1172 2210 1206 2244
rect 1240 2210 1274 2244
rect 1308 2210 1342 2244
rect 1376 2210 1410 2244
rect 1444 2210 1478 2244
rect 1512 2210 1546 2244
rect 84 -90 118 -56
rect 152 -90 186 -56
rect 220 -90 254 -56
rect 288 -90 322 -56
rect 356 -90 390 -56
rect 424 -90 458 -56
rect 492 -90 526 -56
rect 560 -90 594 -56
rect 628 -90 662 -56
rect 696 -90 730 -56
rect 764 -90 798 -56
rect 832 -90 866 -56
rect 900 -90 934 -56
rect 968 -90 1002 -56
rect 1036 -90 1070 -56
rect 1104 -90 1138 -56
rect 1172 -90 1206 -56
rect 1240 -90 1274 -56
rect 1308 -90 1342 -56
rect 1376 -90 1410 -56
rect 1444 -90 1478 -56
rect 1512 -90 1546 -56
<< locali >>
rect -527 2470 2200 2508
rect -527 2368 98 2470
rect 1832 2368 2200 2470
rect -527 2334 2200 2368
rect -527 2117 -286 2334
rect 58 2244 1580 2258
rect 58 2210 78 2244
rect 118 2210 150 2244
rect 186 2210 220 2244
rect 256 2210 288 2244
rect 328 2210 356 2244
rect 400 2210 424 2244
rect 472 2210 492 2244
rect 544 2210 560 2244
rect 616 2210 628 2244
rect 688 2210 696 2244
rect 760 2210 764 2244
rect 866 2210 870 2244
rect 934 2210 942 2244
rect 1002 2210 1014 2244
rect 1070 2210 1086 2244
rect 1138 2210 1158 2244
rect 1206 2210 1230 2244
rect 1274 2210 1302 2244
rect 1342 2210 1374 2244
rect 1410 2210 1444 2244
rect 1480 2210 1512 2244
rect 1552 2210 1580 2244
rect 58 2194 1580 2210
rect -289 111 -286 2117
rect -527 -243 -286 111
rect 1959 1980 2200 2334
rect 2197 -26 2200 1980
rect 58 -56 1580 -42
rect 58 -90 78 -56
rect 118 -90 150 -56
rect 186 -90 220 -56
rect 256 -90 288 -56
rect 328 -90 356 -56
rect 400 -90 424 -56
rect 472 -90 492 -56
rect 544 -90 560 -56
rect 616 -90 628 -56
rect 688 -90 696 -56
rect 760 -90 764 -56
rect 866 -90 870 -56
rect 934 -90 942 -56
rect 1002 -90 1014 -56
rect 1070 -90 1086 -56
rect 1138 -90 1158 -56
rect 1206 -90 1230 -56
rect 1274 -90 1302 -56
rect 1342 -90 1374 -56
rect 1410 -90 1444 -56
rect 1480 -90 1512 -56
rect 1552 -90 1580 -56
rect 58 -106 1580 -90
rect 1959 -243 2200 -26
rect -527 -277 2200 -243
rect -527 -379 41 -277
rect 1775 -379 2200 -277
rect -527 -413 2200 -379
rect -527 -415 -286 -413
<< viali >>
rect 78 2210 84 2244
rect 84 2210 112 2244
rect 150 2210 152 2244
rect 152 2210 184 2244
rect 222 2210 254 2244
rect 254 2210 256 2244
rect 294 2210 322 2244
rect 322 2210 328 2244
rect 366 2210 390 2244
rect 390 2210 400 2244
rect 438 2210 458 2244
rect 458 2210 472 2244
rect 510 2210 526 2244
rect 526 2210 544 2244
rect 582 2210 594 2244
rect 594 2210 616 2244
rect 654 2210 662 2244
rect 662 2210 688 2244
rect 726 2210 730 2244
rect 730 2210 760 2244
rect 798 2210 832 2244
rect 870 2210 900 2244
rect 900 2210 904 2244
rect 942 2210 968 2244
rect 968 2210 976 2244
rect 1014 2210 1036 2244
rect 1036 2210 1048 2244
rect 1086 2210 1104 2244
rect 1104 2210 1120 2244
rect 1158 2210 1172 2244
rect 1172 2210 1192 2244
rect 1230 2210 1240 2244
rect 1240 2210 1264 2244
rect 1302 2210 1308 2244
rect 1308 2210 1336 2244
rect 1374 2210 1376 2244
rect 1376 2210 1408 2244
rect 1446 2210 1478 2244
rect 1478 2210 1480 2244
rect 1518 2210 1546 2244
rect 1546 2210 1552 2244
rect -499 1148 -321 1326
rect 1990 1147 2168 1325
rect 78 -90 84 -56
rect 84 -90 112 -56
rect 150 -90 152 -56
rect 152 -90 184 -56
rect 222 -90 254 -56
rect 254 -90 256 -56
rect 294 -90 322 -56
rect 322 -90 328 -56
rect 366 -90 390 -56
rect 390 -90 400 -56
rect 438 -90 458 -56
rect 458 -90 472 -56
rect 510 -90 526 -56
rect 526 -90 544 -56
rect 582 -90 594 -56
rect 594 -90 616 -56
rect 654 -90 662 -56
rect 662 -90 688 -56
rect 726 -90 730 -56
rect 730 -90 760 -56
rect 798 -90 832 -56
rect 870 -90 900 -56
rect 900 -90 904 -56
rect 942 -90 968 -56
rect 968 -90 976 -56
rect 1014 -90 1036 -56
rect 1036 -90 1048 -56
rect 1086 -90 1104 -56
rect 1104 -90 1120 -56
rect 1158 -90 1172 -56
rect 1172 -90 1192 -56
rect 1230 -90 1240 -56
rect 1240 -90 1264 -56
rect 1302 -90 1308 -56
rect 1308 -90 1336 -56
rect 1374 -90 1376 -56
rect 1376 -90 1408 -56
rect 1446 -90 1478 -56
rect 1478 -90 1480 -56
rect 1518 -90 1546 -56
rect 1546 -90 1552 -56
<< metal1 >>
rect -154 2244 1786 2258
rect -154 2210 78 2244
rect 112 2210 150 2244
rect 184 2210 222 2244
rect 256 2210 294 2244
rect 328 2210 366 2244
rect 400 2210 438 2244
rect 472 2210 510 2244
rect 544 2210 582 2244
rect 616 2210 654 2244
rect 688 2210 726 2244
rect 760 2210 798 2244
rect 832 2210 870 2244
rect 904 2210 942 2244
rect 976 2210 1014 2244
rect 1048 2210 1086 2244
rect 1120 2210 1158 2244
rect 1192 2210 1230 2244
rect 1264 2210 1302 2244
rect 1336 2210 1374 2244
rect 1408 2210 1446 2244
rect 1480 2210 1518 2244
rect 1552 2210 1786 2244
rect -154 2194 1786 2210
rect -154 2081 -62 2194
rect -154 2029 -134 2081
rect -82 2029 -62 2081
rect -154 2017 -62 2029
rect -154 1965 -134 2017
rect -82 1965 -62 2017
rect -527 1327 -286 1373
rect -527 1147 -500 1327
rect -320 1147 -286 1327
rect -527 1103 -286 1147
rect -154 -42 -62 1965
rect 945 2079 1009 2103
rect 945 2027 951 2079
rect 1003 2027 1009 2079
rect 945 2015 1009 2027
rect 945 1963 951 2015
rect 1003 1963 1009 2015
rect 945 1940 1009 1963
rect 1694 2073 1786 2194
rect 1694 2021 1712 2073
rect 1764 2021 1786 2073
rect 1694 2009 1786 2021
rect 1694 1957 1712 2009
rect 1764 1957 1786 2009
rect 313 1755 377 1770
rect 313 1703 319 1755
rect 371 1703 377 1755
rect 313 1691 377 1703
rect 313 1639 319 1691
rect 371 1639 377 1691
rect 313 1627 377 1639
rect 313 1575 319 1627
rect 371 1575 377 1627
rect 313 1560 377 1575
rect 155 1359 219 1373
rect 155 1307 161 1359
rect 213 1307 219 1359
rect 155 1295 219 1307
rect 155 1243 161 1295
rect 213 1243 219 1295
rect 155 1231 219 1243
rect 155 1179 161 1231
rect 213 1179 219 1231
rect 155 1167 219 1179
rect 155 1115 161 1167
rect 213 1115 219 1167
rect 155 1102 219 1115
rect 471 1359 535 1373
rect 471 1307 477 1359
rect 529 1307 535 1359
rect 471 1295 535 1307
rect 471 1243 477 1295
rect 529 1243 535 1295
rect 471 1231 535 1243
rect 471 1179 477 1231
rect 529 1179 535 1231
rect 471 1167 535 1179
rect 471 1115 477 1167
rect 529 1115 535 1167
rect 471 1102 535 1115
rect 787 1359 851 1373
rect 787 1307 793 1359
rect 845 1307 851 1359
rect 787 1295 851 1307
rect 787 1243 793 1295
rect 845 1243 851 1295
rect 787 1231 851 1243
rect 787 1179 793 1231
rect 845 1179 851 1231
rect 787 1167 851 1179
rect 787 1115 793 1167
rect 845 1115 851 1167
rect 787 1102 851 1115
rect 1103 1359 1167 1373
rect 1103 1307 1109 1359
rect 1161 1307 1167 1359
rect 1103 1295 1167 1307
rect 1103 1243 1109 1295
rect 1161 1243 1167 1295
rect 1103 1231 1167 1243
rect 1103 1179 1109 1231
rect 1161 1179 1167 1231
rect 1103 1167 1167 1179
rect 1103 1115 1109 1167
rect 1161 1115 1167 1167
rect 1103 1102 1167 1115
rect 1419 1359 1483 1373
rect 1419 1307 1425 1359
rect 1477 1307 1483 1359
rect 1419 1295 1483 1307
rect 1419 1243 1425 1295
rect 1477 1243 1483 1295
rect 1419 1231 1483 1243
rect 1419 1179 1425 1231
rect 1477 1179 1483 1231
rect 1419 1167 1483 1179
rect 1419 1115 1425 1167
rect 1477 1115 1483 1167
rect 1419 1102 1483 1115
rect -3 256 61 282
rect -3 204 3 256
rect 55 204 61 256
rect -3 192 61 204
rect -3 140 3 192
rect 55 140 61 192
rect -3 115 61 140
rect 629 256 693 282
rect 629 204 635 256
rect 687 204 693 256
rect 629 192 693 204
rect 629 140 635 192
rect 687 140 693 192
rect 629 115 693 140
rect 1261 256 1325 282
rect 1261 204 1267 256
rect 1319 204 1325 256
rect 1261 192 1325 204
rect 1261 140 1267 192
rect 1319 140 1325 192
rect 1261 115 1325 140
rect 1577 256 1641 282
rect 1577 204 1583 256
rect 1635 204 1641 256
rect 1577 192 1641 204
rect 1577 140 1583 192
rect 1635 140 1641 192
rect 1577 115 1641 140
rect 1694 -42 1786 1957
rect 1959 1326 2200 1373
rect 1959 1146 1989 1326
rect 2169 1146 2200 1326
rect 1959 1103 2200 1146
rect -154 -56 1786 -42
rect -154 -90 78 -56
rect 112 -90 150 -56
rect 184 -90 222 -56
rect 256 -90 294 -56
rect 328 -90 366 -56
rect 400 -90 438 -56
rect 472 -90 510 -56
rect 544 -90 582 -56
rect 616 -90 654 -56
rect 688 -90 726 -56
rect 760 -90 798 -56
rect 832 -90 870 -56
rect 904 -90 942 -56
rect 976 -90 1014 -56
rect 1048 -90 1086 -56
rect 1120 -90 1158 -56
rect 1192 -90 1230 -56
rect 1264 -90 1302 -56
rect 1336 -90 1374 -56
rect 1408 -90 1446 -56
rect 1480 -90 1518 -56
rect 1552 -90 1786 -56
rect -154 -106 1786 -90
<< via1 >>
rect -134 2029 -82 2081
rect -134 1965 -82 2017
rect -500 1326 -320 1327
rect -500 1148 -499 1326
rect -499 1148 -321 1326
rect -321 1148 -320 1326
rect -500 1147 -320 1148
rect 951 2027 1003 2079
rect 951 1963 1003 2015
rect 1712 2021 1764 2073
rect 1712 1957 1764 2009
rect 319 1703 371 1755
rect 319 1639 371 1691
rect 319 1575 371 1627
rect 161 1307 213 1359
rect 161 1243 213 1295
rect 161 1179 213 1231
rect 161 1115 213 1167
rect 477 1307 529 1359
rect 477 1243 529 1295
rect 477 1179 529 1231
rect 477 1115 529 1167
rect 793 1307 845 1359
rect 793 1243 845 1295
rect 793 1179 845 1231
rect 793 1115 845 1167
rect 1109 1307 1161 1359
rect 1109 1243 1161 1295
rect 1109 1179 1161 1231
rect 1109 1115 1161 1167
rect 1425 1307 1477 1359
rect 1425 1243 1477 1295
rect 1425 1179 1477 1231
rect 1425 1115 1477 1167
rect 3 204 55 256
rect 3 140 55 192
rect 635 204 687 256
rect 635 140 687 192
rect 1267 204 1319 256
rect 1267 140 1319 192
rect 1583 204 1635 256
rect 1583 140 1635 192
rect 1989 1325 2169 1326
rect 1989 1147 1990 1325
rect 1990 1147 2168 1325
rect 2168 1147 2169 1325
rect 1989 1146 2169 1147
<< metal2 >>
rect -154 2081 1786 2104
rect -154 2029 -134 2081
rect -82 2079 1786 2081
rect -82 2029 951 2079
rect -154 2027 951 2029
rect 1003 2073 1786 2079
rect 1003 2027 1712 2073
rect -154 2021 1712 2027
rect 1764 2021 1786 2073
rect -154 2017 1786 2021
rect -154 1965 -134 2017
rect -82 2015 1786 2017
rect -82 1965 951 2015
rect -154 1963 951 1965
rect 1003 2009 1786 2015
rect 1003 1963 1712 2009
rect -154 1957 1712 1963
rect 1764 1957 1786 2009
rect -154 1938 1786 1957
rect 0 1755 1638 1772
rect 0 1703 319 1755
rect 371 1703 1638 1755
rect 0 1691 1638 1703
rect 0 1639 319 1691
rect 371 1639 1638 1691
rect 0 1627 1638 1639
rect 0 1575 319 1627
rect 371 1575 1638 1627
rect 0 1556 1638 1575
rect -527 1359 2200 1373
rect -527 1327 161 1359
rect -527 1147 -500 1327
rect -320 1307 161 1327
rect 213 1307 477 1359
rect 529 1307 793 1359
rect 845 1307 1109 1359
rect 1161 1307 1425 1359
rect 1477 1326 2200 1359
rect 1477 1307 1989 1326
rect -320 1295 1989 1307
rect -320 1243 161 1295
rect 213 1243 477 1295
rect 529 1243 793 1295
rect 845 1243 1109 1295
rect 1161 1243 1425 1295
rect 1477 1243 1989 1295
rect -320 1231 1989 1243
rect -320 1179 161 1231
rect 213 1179 477 1231
rect 529 1179 793 1231
rect 845 1179 1109 1231
rect 1161 1179 1425 1231
rect 1477 1179 1989 1231
rect -320 1167 1989 1179
rect -320 1147 161 1167
rect -527 1115 161 1147
rect 213 1115 477 1167
rect 529 1115 793 1167
rect 845 1115 1109 1167
rect 1161 1115 1425 1167
rect 1477 1146 1989 1167
rect 2169 1146 2200 1326
rect 1477 1115 2200 1146
rect -527 1103 2200 1115
rect -3 256 1641 282
rect -3 204 3 256
rect 55 204 635 256
rect 687 204 1267 256
rect 1319 204 1583 256
rect 1635 204 1641 256
rect -3 192 1641 204
rect -3 140 3 192
rect 55 140 635 192
rect 687 140 1267 192
rect 1319 140 1583 192
rect 1635 140 1641 192
rect -3 116 1641 140
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_0
timestamp 1667803582
transform 1 0 1530 0 1 1076
box -134 -1076 134 1076
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_1
timestamp 1667803582
transform 1 0 1214 0 1 1076
box -134 -1076 134 1076
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_2
timestamp 1667803582
transform 1 0 1372 0 1 1076
box -134 -1076 134 1076
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_3
timestamp 1667803582
transform 1 0 1056 0 1 1076
box -134 -1076 134 1076
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_4
timestamp 1667803582
transform 1 0 740 0 1 1076
box -134 -1076 134 1076
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_5
timestamp 1667803582
transform 1 0 898 0 1 1076
box -134 -1076 134 1076
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_6
timestamp 1667803582
transform 1 0 424 0 1 1076
box -134 -1076 134 1076
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_7
timestamp 1667803582
transform 1 0 582 0 1 1076
box -134 -1076 134 1076
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_8
timestamp 1667803582
transform 1 0 108 0 1 1076
box -134 -1076 134 1076
use sky130_fd_pr__nfet_01v8_RC9KLY  sky130_fd_pr__nfet_01v8_RC9KLY_9
timestamp 1667803582
transform 1 0 266 0 1 1076
box -134 -1076 134 1076
<< labels >>
flabel metal2 s 108 177 108 177 0 FreeSans 1250 0 0 0 D3
port 1 nsew
flabel metal2 s 88 1226 88 1226 0 FreeSans 1250 0 0 0 S
port 2 nsew
flabel metal2 s 262 2027 262 2027 0 FreeSans 1250 0 0 0 D1
port 3 nsew
flabel metal2 s 266 1667 266 1667 0 FreeSans 1250 0 0 0 D2
port 4 nsew
<< end >>
