magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< nwell >>
rect -121 1057 898 1162
rect -135 937 898 1057
rect -472 343 898 937
rect -662 38 898 343
rect -655 0 802 38
<< poly >>
rect 96 1119 434 1197
rect 482 1126 818 1197
rect 291 1100 317 1119
rect 80 2 416 75
rect 464 2 801 74
rect 98 -44 416 2
rect 482 -44 801 2
rect 98 -110 434 -44
rect 482 -110 818 -44
rect 80 -720 416 -653
rect 464 -720 800 -654
<< viali >>
rect -528 46 -494 80
<< metal1 >>
rect -65 1141 434 1188
rect 560 1141 977 1187
rect -2581 235 -247 331
rect -554 162 -470 175
rect -554 110 -539 162
rect -487 110 -470 162
rect -554 80 -470 110
rect -554 46 -528 80
rect -494 46 -470 80
rect -554 31 -470 46
rect -65 59 -19 1141
rect 117 1073 202 1100
rect 117 1021 134 1073
rect 186 1021 202 1073
rect 117 1009 202 1021
rect 117 957 134 1009
rect 186 957 202 1009
rect 117 923 202 957
rect 310 1069 395 1100
rect 310 1017 327 1069
rect 379 1017 395 1069
rect 310 1005 395 1017
rect 310 953 327 1005
rect 379 953 395 1005
rect 310 924 395 953
rect 507 866 580 902
rect 507 814 516 866
rect 568 814 580 866
rect 507 780 580 814
rect 700 867 782 902
rect 700 815 715 867
rect 767 815 782 867
rect 700 780 782 815
rect 41 381 107 396
rect 41 329 48 381
rect 100 329 107 381
rect 41 309 107 329
rect 213 380 298 396
rect 213 328 231 380
rect 283 328 298 380
rect 213 309 298 328
rect 416 377 483 395
rect 416 325 420 377
rect 472 325 483 377
rect 416 309 483 325
rect 608 378 674 395
rect 608 326 614 378
rect 666 326 674 378
rect 608 309 674 326
rect 793 378 862 396
rect 793 326 801 378
rect 853 326 862 378
rect 793 309 862 326
rect 931 59 977 1141
rect -65 0 338 59
rect 468 35 977 59
rect 468 13 602 35
rect -2289 -47 -2138 0
rect -724 -54 338 0
rect 560 -17 602 13
rect 654 -17 977 35
rect -724 -83 434 -54
rect -65 -100 434 -83
rect 560 -100 977 -17
rect -2581 -309 -247 -213
rect -65 -664 -19 -100
rect 34 -171 100 -147
rect 34 -223 41 -171
rect 93 -223 100 -171
rect 34 -235 100 -223
rect 34 -287 41 -235
rect 93 -287 100 -235
rect 34 -309 100 -287
rect 218 -171 293 -147
rect 218 -223 228 -171
rect 280 -223 293 -171
rect 218 -235 293 -223
rect 218 -287 228 -235
rect 280 -287 293 -235
rect 218 -308 293 -287
rect 412 -171 484 -147
rect 412 -223 417 -171
rect 469 -223 484 -171
rect 412 -235 484 -223
rect 412 -287 417 -235
rect 469 -287 484 -235
rect 412 -309 484 -287
rect 607 -171 677 -147
rect 607 -223 614 -171
rect 666 -223 677 -171
rect 607 -235 677 -223
rect 607 -287 614 -235
rect 666 -287 677 -235
rect 607 -309 677 -287
rect 800 -171 862 -147
rect 800 -223 807 -171
rect 859 -223 862 -171
rect 800 -235 862 -223
rect 800 -287 807 -235
rect 859 -287 862 -235
rect 800 -309 862 -287
rect 125 -428 195 -387
rect 125 -480 133 -428
rect 185 -480 195 -428
rect 125 -492 195 -480
rect 125 -544 133 -492
rect 185 -544 195 -492
rect 125 -586 195 -544
rect 316 -432 388 -387
rect 316 -484 327 -432
rect 379 -484 388 -432
rect 316 -496 388 -484
rect 316 -548 327 -496
rect 379 -548 388 -496
rect 316 -588 388 -548
rect 505 -429 580 -387
rect 505 -481 516 -429
rect 568 -481 580 -429
rect 505 -493 580 -481
rect 505 -545 516 -493
rect 568 -545 580 -493
rect 505 -587 580 -545
rect 698 -398 769 -387
rect 698 -450 707 -398
rect 759 -450 769 -398
rect 698 -462 769 -450
rect 698 -514 707 -462
rect 759 -514 769 -462
rect 698 -526 769 -514
rect 698 -578 707 -526
rect 759 -578 769 -526
rect 698 -588 769 -578
rect 931 -664 977 -100
rect -65 -710 338 -664
rect 464 -711 977 -664
<< via1 >>
rect -539 110 -487 162
rect 134 1021 186 1073
rect 134 957 186 1009
rect 327 1017 379 1069
rect 327 953 379 1005
rect 516 814 568 866
rect 715 815 767 867
rect 48 329 100 381
rect 231 328 283 380
rect 420 325 472 377
rect 614 326 666 378
rect 801 326 853 378
rect 602 -17 654 35
rect 41 -223 93 -171
rect 41 -287 93 -235
rect 228 -223 280 -171
rect 228 -287 280 -235
rect 417 -223 469 -171
rect 417 -287 469 -235
rect 614 -223 666 -171
rect 614 -287 666 -235
rect 807 -223 859 -171
rect 807 -287 859 -235
rect 133 -480 185 -428
rect 133 -544 185 -492
rect 327 -484 379 -432
rect 327 -548 379 -496
rect 516 -481 568 -429
rect 516 -545 568 -493
rect 707 -450 759 -398
rect 707 -514 759 -462
rect 707 -578 759 -526
<< metal2 >>
rect 118 1073 977 1100
rect 118 1021 134 1073
rect 186 1069 977 1073
rect 186 1021 327 1069
rect 118 1017 327 1021
rect 379 1017 977 1069
rect 118 1009 977 1017
rect 118 957 134 1009
rect 186 1005 977 1009
rect 186 957 327 1005
rect 118 953 327 957
rect 379 953 977 1005
rect 118 940 977 953
rect 118 923 400 940
rect 507 888 782 902
rect -67 867 782 888
rect -67 866 715 867
rect -67 814 516 866
rect 568 815 715 866
rect 767 815 782 867
rect 568 814 782 815
rect -67 780 782 814
rect -67 375 -13 780
rect -87 368 -13 375
rect -87 312 -77 368
rect -21 312 -13 368
rect -87 303 -13 312
rect 42 381 862 396
rect 42 329 48 381
rect 100 380 862 381
rect 100 329 231 380
rect 42 328 231 329
rect 283 378 862 380
rect 283 377 614 378
rect 283 328 420 377
rect 42 325 420 328
rect 472 326 614 377
rect 666 326 801 378
rect 853 326 862 378
rect 472 325 862 326
rect 42 309 862 325
rect -554 162 675 228
rect -554 110 -539 162
rect -487 118 675 162
rect -487 110 -470 118
rect -554 31 -470 110
rect -87 51 -13 61
rect -87 -5 -78 51
rect -22 -5 -13 51
rect -87 -14 -13 -5
rect -67 -388 -13 -14
rect 581 35 675 118
rect 581 -17 602 35
rect 654 -17 675 35
rect 581 -40 675 -17
rect 754 -147 862 309
rect 34 -171 862 -147
rect 34 -223 41 -171
rect 93 -223 228 -171
rect 280 -223 417 -171
rect 469 -223 614 -171
rect 666 -223 807 -171
rect 859 -223 862 -171
rect 34 -235 862 -223
rect 34 -287 41 -235
rect 93 -287 228 -235
rect 280 -287 417 -235
rect 469 -287 614 -235
rect 666 -287 807 -235
rect 859 -287 862 -235
rect 34 -309 862 -287
rect 927 -387 977 940
rect 125 -388 387 -387
rect -67 -428 387 -388
rect -67 -480 133 -428
rect 185 -432 387 -428
rect 185 -480 327 -432
rect -67 -484 327 -480
rect 379 -484 387 -432
rect -67 -492 387 -484
rect -67 -544 133 -492
rect 185 -496 387 -492
rect 185 -544 327 -496
rect -67 -548 327 -544
rect 379 -548 387 -496
rect -67 -587 387 -548
rect 501 -398 977 -387
rect 501 -429 707 -398
rect 501 -481 516 -429
rect 568 -450 707 -429
rect 759 -450 977 -398
rect 568 -462 977 -450
rect 568 -481 707 -462
rect 501 -493 707 -481
rect 501 -545 516 -493
rect 568 -514 707 -493
rect 759 -514 977 -462
rect 568 -526 977 -514
rect 568 -545 707 -526
rect 501 -578 707 -545
rect 759 -578 977 -526
rect 501 -587 977 -578
<< via2 >>
rect -77 312 -21 368
rect -78 -5 -22 51
<< metal3 >>
rect -87 368 -13 375
rect -87 312 -77 368
rect -21 312 -13 368
rect -87 51 -13 312
rect -87 -5 -78 51
rect -22 -5 -13 51
rect -87 -14 -13 -5
use sky130_fd_pr__nfet_01v8_WWN8PW  sky130_fd_pr__nfet_01v8_WWN8PW_0
timestamp 1667803582
transform 1 0 641 0 1 -382
box -247 -338 247 338
use sky130_fd_pr__nfet_01v8_WWN8PW  sky130_fd_pr__nfet_01v8_WWN8PW_1
timestamp 1667803582
transform 1 0 257 0 1 -382
box -247 -338 247 338
use sky130_fd_pr__pfet_01v8_52DJHB  sky130_fd_pr__pfet_01v8_52DJHB_0
timestamp 1667803582
transform 1 0 641 0 1 600
box -257 -600 257 600
use sky130_fd_pr__pfet_01v8_52DJHB  sky130_fd_pr__pfet_01v8_52DJHB_1
timestamp 1667803582
transform 1 0 257 0 1 600
box -257 -600 257 600
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0
timestamp 1667803582
transform 1 0 -2581 0 1 -261
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1667803582
transform 1 0 -339 0 1 -261
box -38 -48 130 592
<< labels >>
flabel metal2 s 159 1006 159 1006 0 FreeSans 600 0 0 0 VREF_P
port 1 nsew
flabel metal2 s 546 865 546 865 0 FreeSans 600 0 0 0 VREF_N
port 2 nsew
flabel metal2 s 260 363 260 363 0 FreeSans 600 0 0 0 VOUT
port 3 nsew
flabel metal1 s -1590 282 -1590 282 0 FreeSans 800 0 0 0 VDD
port 4 nsew
flabel metal1 s -1671 -271 -1671 -271 0 FreeSans 800 0 0 0 VSS
port 5 nsew
flabel metal1 s -2230 -19 -2230 -19 0 FreeSans 800 0 0 0 VIN
port 6 nsew
<< end >>
