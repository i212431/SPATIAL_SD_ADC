magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< locali >>
rect 1815 1294 1953 1325
<< metal1 >>
rect 187 2445 640 2491
rect 42 2381 105 2410
rect 42 2329 48 2381
rect 100 2329 105 2381
rect 42 2317 105 2329
rect 42 2265 48 2317
rect 100 2265 105 2317
rect 42 2236 105 2265
rect 230 2381 299 2410
rect 230 2329 238 2381
rect 290 2329 299 2381
rect 230 2317 299 2329
rect 230 2265 238 2317
rect 290 2265 299 2317
rect 230 2235 299 2265
rect 422 2380 491 2412
rect 422 2328 431 2380
rect 483 2328 491 2380
rect 422 2316 491 2328
rect 422 2264 431 2316
rect 483 2264 491 2316
rect 422 2236 491 2264
rect 134 2053 201 2078
rect 134 2001 142 2053
rect 194 2001 201 2053
rect 134 1989 201 2001
rect 134 1937 142 1989
rect 194 1937 201 1989
rect 134 1912 201 1937
rect 327 2053 394 2078
rect 327 2001 335 2053
rect 387 2001 394 2053
rect 327 1989 394 2001
rect 327 1937 335 1989
rect 387 1937 394 1989
rect 327 1912 394 1937
rect 594 1880 640 2445
rect 1828 2443 2277 2488
rect 1684 2381 1751 2410
rect 1684 2329 1691 2381
rect 1743 2329 1751 2381
rect 1684 2317 1751 2329
rect 1684 2265 1691 2317
rect 1743 2265 1751 2317
rect 1684 2236 1751 2265
rect 1877 2382 1944 2411
rect 1877 2330 1885 2382
rect 1937 2330 1944 2382
rect 1877 2318 1944 2330
rect 1877 2266 1885 2318
rect 1937 2266 1944 2318
rect 1877 2235 1944 2266
rect 2069 2382 2133 2410
rect 2069 2330 2075 2382
rect 2127 2330 2133 2382
rect 2069 2318 2133 2330
rect 2069 2266 2075 2318
rect 2127 2266 2133 2318
rect 2069 2236 2133 2266
rect 1779 2135 1848 2154
rect 1779 2083 1786 2135
rect 1838 2083 1848 2135
rect 1779 2071 1848 2083
rect 1779 2019 1786 2071
rect 1838 2019 1848 2071
rect 1779 2007 1848 2019
rect 1779 1955 1786 2007
rect 1838 1955 1848 2007
rect 1779 1937 1848 1955
rect 1972 2136 2042 2155
rect 1972 2084 1980 2136
rect 2032 2084 2042 2136
rect 1972 2072 2042 2084
rect 1972 2020 1980 2072
rect 2032 2020 2042 2072
rect 1972 2008 2042 2020
rect 1972 1956 1980 2008
rect 2032 1956 2042 2008
rect 1972 1936 2042 1956
rect 87 1872 640 1880
rect 2232 1876 2277 2443
rect 87 1834 290 1872
rect 277 1820 290 1834
rect 342 1820 354 1872
rect 406 1820 418 1872
rect 470 1834 640 1872
rect 1733 1860 2277 1876
rect 470 1820 483 1834
rect 1733 1831 1835 1860
rect 277 1803 483 1820
rect 1800 1808 1835 1831
rect 1887 1808 1899 1860
rect 1951 1831 2277 1860
rect 1951 1808 1988 1831
rect 1800 1794 1988 1808
rect -110 1572 2246 1594
rect -110 1520 1315 1572
rect 1367 1520 1379 1572
rect 1431 1520 2246 1572
rect -110 1498 2246 1520
rect 1802 1371 2183 1373
rect 1801 1348 2183 1371
rect 1801 1296 1838 1348
rect 1890 1296 1902 1348
rect 1954 1296 2183 1348
rect 1801 1283 2183 1296
rect 1801 1281 1989 1283
rect -441 1251 201 1254
rect -441 1225 206 1251
rect 150 1091 206 1225
rect -110 954 2394 1050
rect 105 703 481 720
rect 1823 711 2045 719
rect 105 651 324 703
rect 376 651 388 703
rect 440 651 481 703
rect 105 634 481 651
rect 1822 699 2047 711
rect 1822 647 1843 699
rect 1895 647 1907 699
rect 1959 647 1971 699
rect 2023 647 2047 699
rect 1822 637 2047 647
rect 38 482 2394 506
rect 38 430 1317 482
rect 1369 430 1381 482
rect 1433 430 2394 482
rect 38 410 2394 430
<< via1 >>
rect 48 2329 100 2381
rect 48 2265 100 2317
rect 238 2329 290 2381
rect 238 2265 290 2317
rect 431 2328 483 2380
rect 431 2264 483 2316
rect 142 2001 194 2053
rect 142 1937 194 1989
rect 335 2001 387 2053
rect 335 1937 387 1989
rect 1691 2329 1743 2381
rect 1691 2265 1743 2317
rect 1885 2330 1937 2382
rect 1885 2266 1937 2318
rect 2075 2330 2127 2382
rect 2075 2266 2127 2318
rect 1786 2083 1838 2135
rect 1786 2019 1838 2071
rect 1786 1955 1838 2007
rect 1980 2084 2032 2136
rect 1980 2020 2032 2072
rect 1980 1956 2032 2008
rect 290 1820 342 1872
rect 354 1820 406 1872
rect 418 1820 470 1872
rect 1835 1808 1887 1860
rect 1899 1808 1951 1860
rect 1315 1520 1367 1572
rect 1379 1520 1431 1572
rect 1838 1296 1890 1348
rect 1902 1296 1954 1348
rect 324 651 376 703
rect 388 651 440 703
rect 1843 647 1895 699
rect 1907 647 1959 699
rect 1971 647 2023 699
rect 1317 430 1369 482
rect 1381 430 1433 482
<< metal2 >>
rect 422 2411 491 2412
rect 49 2410 491 2411
rect 42 2382 2133 2410
rect 42 2381 1885 2382
rect 42 2329 48 2381
rect 100 2329 238 2381
rect 290 2380 1691 2381
rect 290 2329 431 2380
rect 42 2328 431 2329
rect 483 2329 1691 2380
rect 1743 2330 1885 2381
rect 1937 2330 2075 2382
rect 2127 2330 2133 2382
rect 1743 2329 2133 2330
rect 483 2328 2133 2329
rect 42 2318 2133 2328
rect 42 2317 1885 2318
rect 42 2265 48 2317
rect 100 2265 238 2317
rect 290 2316 1691 2317
rect 290 2265 431 2316
rect 42 2264 431 2265
rect 483 2265 1691 2316
rect 1743 2266 1885 2317
rect 1937 2266 2075 2318
rect 2127 2266 2133 2318
rect 1743 2265 2133 2266
rect 483 2264 2133 2265
rect 42 2236 2133 2264
rect 1687 2136 2480 2155
rect 1687 2135 1980 2136
rect 1687 2083 1786 2135
rect 1838 2084 1980 2135
rect 2032 2084 2480 2136
rect 1838 2083 2480 2084
rect -231 2053 480 2078
rect -231 2001 142 2053
rect 194 2001 335 2053
rect 387 2001 480 2053
rect -231 1989 480 2001
rect -231 1937 142 1989
rect 194 1937 335 1989
rect 387 1937 480 1989
rect -231 1912 480 1937
rect 1687 2072 2480 2083
rect 1687 2071 1980 2072
rect 1687 2019 1786 2071
rect 1838 2020 1980 2071
rect 2032 2020 2480 2072
rect 1838 2019 2480 2020
rect 1687 2008 2480 2019
rect 1687 2007 1980 2008
rect 1687 1955 1786 2007
rect 1838 1956 1980 2007
rect 2032 1956 2480 2008
rect 1838 1955 2480 1956
rect 1687 1936 2480 1955
rect -231 1874 -65 1912
rect -397 1708 -65 1874
rect 277 1872 483 1880
rect 1802 1874 1989 1888
rect 277 1820 290 1872
rect 342 1820 354 1872
rect 406 1820 418 1872
rect 470 1820 483 1872
rect 277 1803 483 1820
rect -689 1343 -505 1364
rect -689 1287 -665 1343
rect -609 1287 -585 1343
rect -529 1287 -505 1343
rect -689 1266 -505 1287
rect 278 703 483 1803
rect 1800 1860 1989 1874
rect 1800 1808 1835 1860
rect 1887 1808 1899 1860
rect 1951 1808 1989 1860
rect 1800 1794 1989 1808
rect 278 651 324 703
rect 376 651 388 703
rect 440 651 483 703
rect 278 636 483 651
rect 1284 1572 1465 1594
rect 1284 1520 1315 1572
rect 1367 1520 1379 1572
rect 1431 1520 1465 1572
rect 1284 482 1465 1520
rect 1802 1373 1989 1794
rect 1802 1348 2183 1373
rect 1802 1296 1838 1348
rect 1890 1296 1902 1348
rect 1954 1296 2183 1348
rect 1802 1283 2183 1296
rect 2261 1080 2480 1936
rect 2261 861 2992 1080
rect 1823 699 2182 713
rect 1823 647 1843 699
rect 1895 647 1907 699
rect 1959 647 1971 699
rect 2023 647 2182 699
rect 1823 635 2182 647
rect 3023 618 3248 781
rect 1284 430 1317 482
rect 1369 430 1381 482
rect 1433 430 1465 482
rect 1284 410 1465 430
rect 2795 550 2973 551
rect 2795 414 2816 550
rect 2952 414 2973 550
rect -1033 376 -738 395
rect -1033 240 -1015 376
rect -879 368 -738 376
rect -879 336 -695 368
rect -879 280 -834 336
rect -778 280 -754 336
rect -698 280 -695 336
rect -879 248 -695 280
rect -879 240 -738 248
rect -1033 223 -738 240
<< via2 >>
rect -665 1287 -609 1343
rect -585 1287 -529 1343
rect 2816 414 2952 550
rect -1015 240 -879 376
rect -834 280 -778 336
rect -754 280 -698 336
<< metal3 >>
rect -705 1343 -493 1378
rect -705 1287 -665 1343
rect -609 1287 -585 1343
rect -529 1287 -493 1343
rect -705 1251 -493 1287
rect 2784 550 3441 570
rect 2784 414 2816 550
rect 2952 517 3441 550
rect 2952 453 3327 517
rect 3391 453 3441 517
rect 2952 414 3441 453
rect -936 394 -673 395
rect 2784 394 3441 414
rect -1032 380 -673 394
rect -1032 236 -1018 380
rect -874 336 -673 380
rect -874 280 -834 336
rect -778 280 -754 336
rect -698 280 -673 336
rect -874 236 -673 280
rect -1032 224 -673 236
rect -936 223 -673 224
<< via3 >>
rect 3327 453 3391 517
rect -1018 376 -874 380
rect -1018 240 -1015 376
rect -1015 240 -879 376
rect -879 240 -874 376
rect -1018 236 -874 240
<< metal4 >>
rect 3277 517 4205 570
rect 3277 453 3327 517
rect 3391 453 4205 517
rect -1032 380 -863 394
rect 3277 380 4205 453
rect -1032 236 -1018 380
rect -874 236 -863 380
rect -1032 -642 -863 236
rect 4016 -6004 4205 380
use T_Gate  T_Gate_0
timestamp 1667803582
transform -1 0 -358 0 -1 2004
box -2642 0 541 1919
use T_Gate  T_Gate_1
timestamp 1667803582
transform 1 0 2642 0 1 0
box -2642 0 541 1919
use sky130_fd_pr__cap_mim_m3_1_4RKXMF  sky130_fd_pr__cap_mim_m3_1_4RKXMF_0
timestamp 1667803582
transform 1 0 1130 0 1 -3350
box -2950 -2900 2949 2900
use sky130_fd_pr__nfet_01v8_FR7DL7  sky130_fd_pr__nfet_01v8_FR7DL7_0
timestamp 1667803582
transform 1 0 1910 0 1 2160
box -349 -450 349 450
use sky130_fd_pr__nfet_01v8_FR7DL7  sky130_fd_pr__nfet_01v8_FR7DL7_1
timestamp 1667803582
transform 1 0 264 0 1 2162
box -349 -450 349 450
<< labels >>
flabel metal2 s 1361 1548 1361 1548 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal1 s 951 995 951 995 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal2 s 1076 2334 1076 2334 0 FreeSans 2000 0 0 0 VREF
port 3 nsew
flabel metal3 s -589 1313 -589 1313 0 FreeSans 2000 0 0 0 VIN
port 4 nsew
flabel metal2 s 3207 695 3207 695 0 FreeSans 2000 0 0 0 VOUT
port 5 nsew
flabel metal2 s 1887 1832 1887 1832 0 FreeSans 2000 0 0 0 PH1
port 6 nsew
flabel metal2 s 1917 672 1917 672 0 FreeSans 2000 0 0 0 PH2
port 7 nsew
<< end >>
