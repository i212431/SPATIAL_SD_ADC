magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< metal1 >>
rect -4428 11060 -4186 11062
rect -4428 11008 -4397 11060
rect -4345 11008 -4333 11060
rect -4281 11008 -4269 11060
rect -4217 11008 -4186 11060
rect -4428 11006 -4186 11008
<< via1 >>
rect -4397 11008 -4345 11060
rect -4333 11008 -4281 11060
rect -4269 11008 -4217 11060
<< metal2 >>
rect -1714 12439 1388 12443
rect -3149 12265 1388 12439
rect -1714 11502 1388 12265
rect -3853 11461 -3716 11489
rect -3717 11245 -3716 11461
rect -3853 11218 -3716 11245
rect -4539 11145 -4082 11207
rect -4539 10929 -4455 11145
rect -4159 10929 -4082 11145
rect -4539 10881 -4082 10929
rect -1937 10647 330 10808
rect 1045 10798 1771 10830
rect 1045 10342 1060 10798
rect 1756 10342 1771 10798
rect 1045 10310 1771 10342
<< via2 >>
rect -3853 11245 -3717 11461
rect -4455 11060 -4159 11145
rect -4455 11008 -4397 11060
rect -4397 11008 -4345 11060
rect -4345 11008 -4333 11060
rect -4333 11008 -4281 11060
rect -4281 11008 -4269 11060
rect -4269 11008 -4217 11060
rect -4217 11008 -4159 11060
rect -4455 10929 -4159 11008
rect 1060 10342 1756 10798
<< metal3 >>
rect 6451 13452 7361 13487
rect -3874 12768 3528 12970
rect 6451 12828 6474 13452
rect 7338 12828 7361 13452
rect 6451 12793 7361 12828
rect -3874 11461 -3672 12768
rect -3874 11245 -3853 11461
rect -3717 11245 -3672 11461
rect -4539 11149 -4082 11207
rect -3874 11187 -3672 11245
rect -4539 10925 -4459 11149
rect -4155 10925 -4082 11149
rect -4539 10881 -4082 10925
rect 974 10802 1835 10904
rect 974 10338 1056 10802
rect 1760 10338 1835 10802
rect 974 10243 1835 10338
<< via3 >>
rect 6474 12828 7338 13452
rect -4459 11145 -4155 11149
rect -4459 10929 -4455 11145
rect -4455 10929 -4159 11145
rect -4159 10929 -4155 11145
rect -4459 10925 -4155 10929
rect 1056 10798 1760 10802
rect 1056 10342 1060 10798
rect 1060 10342 1756 10798
rect 1756 10342 1760 10798
rect 1056 10338 1760 10342
<< metal4 >>
rect 6303 13452 7475 13621
rect 6303 13347 6474 13452
rect -4544 12885 6474 13347
rect -4544 11174 -4082 12885
rect 6303 12828 6474 12885
rect 7338 12828 7475 13452
rect 6303 12672 7475 12828
rect -4539 11149 -4082 11174
rect -4539 10925 -4459 11149
rect -4155 10925 -4082 11149
rect -4539 10881 -4082 10925
rect 973 10802 1838 10903
rect 973 10338 1056 10802
rect 1760 10338 1838 10802
rect 973 6230 1838 10338
rect 2624 7032 5479 7277
rect 2624 4578 8777 7032
rect 2624 4004 5479 4578
rect 6323 2850 8777 4578
rect 6323 2764 20947 2850
rect 22076 2764 24491 10997
rect 6323 396 24491 2764
rect 18920 349 24491 396
use OpampM  OpampM_0
timestamp 1667803582
transform 1 0 9213 0 1 10004
box -9221 -10004 21004 11474
use co  co_0
timestamp 1667803582
transform 1 0 -5156 0 1 10029
box -1820 -6250 4205 2612
use sky130_fd_pr__cap_mim_m3_1_D7CHNQ  sky130_fd_pr__cap_mim_m3_1_D7CHNQ_0
timestamp 1667803582
transform 1 0 1069 0 1 5648
box -1650 -1600 1649 1600
<< end >>
