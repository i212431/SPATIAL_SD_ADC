magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< locali >>
rect 10 216 24 258
rect 715 215 789 258
rect 1485 215 1562 258
rect 2214 214 2276 258
<< metal1 >>
rect 0 495 2409 592
rect 0 -48 2409 47
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_0
timestamp 1667803582
transform 1 0 1544 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_1
timestamp 1667803582
transform 1 0 0 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_2
timestamp 1667803582
transform 1 0 770 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1667803582
transform 1 0 2317 0 1 0
box -38 -48 130 592
<< labels >>
flabel metal1 s 1070 542 1070 542 0 FreeSans 200 0 0 0 VDD
port 1 nsew
flabel metal1 s 1087 -18 1087 -18 0 FreeSans 200 0 0 0 VSS
port 2 nsew
flabel locali s 2266 234 2266 234 0 FreeSans 1000 0 0 0 VOUT
port 3 nsew
flabel locali s 14 238 14 238 0 FreeSans 1000 0 0 0 VIN
port 4 nsew
<< end >>
