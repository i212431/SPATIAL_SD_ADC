magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< error_p >>
rect -29 141 29 147
rect -29 107 -17 141
rect -29 101 29 107
<< pwell >>
rect -201 -269 201 269
<< nmos >>
rect -15 -131 15 69
<< ndiff >>
rect -73 54 -15 69
rect -73 20 -61 54
rect -27 20 -15 54
rect -73 -14 -15 20
rect -73 -48 -61 -14
rect -27 -48 -15 -14
rect -73 -82 -15 -48
rect -73 -116 -61 -82
rect -27 -116 -15 -82
rect -73 -131 -15 -116
rect 15 54 73 69
rect 15 20 27 54
rect 61 20 73 54
rect 15 -14 73 20
rect 15 -48 27 -14
rect 61 -48 73 -14
rect 15 -82 73 -48
rect 15 -116 27 -82
rect 61 -116 73 -82
rect 15 -131 73 -116
<< ndiffc >>
rect -61 20 -27 54
rect -61 -48 -27 -14
rect -61 -116 -27 -82
rect 27 20 61 54
rect 27 -48 61 -14
rect 27 -116 61 -82
<< psubdiff >>
rect -175 209 175 243
rect -175 -209 -141 209
rect 141 -209 175 209
rect -175 -243 175 -209
<< poly >>
rect -33 141 33 157
rect -33 107 -17 141
rect 17 107 33 141
rect -33 91 33 107
rect -15 69 15 91
rect -15 -157 15 -131
<< polycont >>
rect -17 107 17 141
<< locali >>
rect -175 209 175 243
rect -175 -209 -141 209
rect -33 107 -17 141
rect 17 107 33 141
rect -61 54 -27 73
rect -61 -14 -27 -12
rect -61 -50 -27 -48
rect -61 -135 -27 -116
rect 27 54 61 73
rect 27 -14 61 -12
rect 27 -50 61 -48
rect 27 -135 61 -116
rect 141 -209 175 209
rect -175 -243 175 -209
<< viali >>
rect -17 107 17 141
rect -61 20 -27 22
rect -61 -12 -27 20
rect -61 -82 -27 -50
rect -61 -84 -27 -82
rect 27 20 61 22
rect 27 -12 61 20
rect 27 -82 61 -50
rect 27 -84 61 -82
<< metal1 >>
rect -29 141 29 147
rect -29 107 -17 141
rect 17 107 29 141
rect -29 101 29 107
rect -67 22 -21 69
rect -67 -12 -61 22
rect -27 -12 -21 22
rect -67 -50 -21 -12
rect -67 -84 -61 -50
rect -27 -84 -21 -50
rect -67 -131 -21 -84
rect 21 22 67 69
rect 21 -12 27 22
rect 61 -12 67 22
rect 21 -50 67 -12
rect 21 -84 27 -50
rect 61 -84 67 -50
rect 21 -131 67 -84
<< properties >>
string FIXED_BBOX -158 -226 158 226
<< end >>
