magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< locali >>
rect 2611 1366 2727 1395
rect 2611 1332 2653 1366
rect 2687 1332 2727 1366
rect 2611 1303 2727 1332
rect 2624 878 2664 1303
rect 2624 838 2851 878
rect 5014 835 5303 869
rect 6682 836 6831 875
rect 9086 873 9294 875
rect 9086 854 9349 873
rect 5522 832 5556 833
rect 9086 820 9276 854
rect 9310 820 9349 854
rect 9086 818 9349 820
rect 9244 797 9349 818
rect 9246 790 9349 797
rect 2782 282 2818 306
rect 2852 282 2862 306
rect 5154 282 5391 322
rect 6801 310 6839 311
rect 2782 214 2862 282
rect 6801 276 6803 310
rect 6837 276 6839 310
rect 8014 288 8126 322
rect 8014 282 8150 288
rect 6801 275 6839 276
<< viali >>
rect 2653 1332 2687 1366
rect 5522 798 5556 832
rect 9276 820 9310 854
rect 2818 282 2852 316
rect 5114 288 5148 322
rect 6803 276 6837 310
rect 7978 282 8012 316
rect 8126 288 8160 322
rect 10423 282 10457 316
<< metal1 >>
rect 2611 1375 2727 1395
rect 2611 1323 2643 1375
rect 2695 1323 2727 1375
rect 2611 1303 2727 1323
rect 2353 1212 2894 1250
rect 2353 1194 11505 1212
rect 2350 1191 11505 1194
rect 2350 1189 10869 1191
rect 2350 1137 8279 1189
rect 8331 1137 8343 1189
rect 8395 1137 8407 1189
rect 8459 1137 8471 1189
rect 8523 1137 8535 1189
rect 8587 1137 8599 1189
rect 8651 1139 10869 1189
rect 10921 1139 10933 1191
rect 10985 1139 10997 1191
rect 11049 1139 11505 1191
rect 8651 1137 11505 1139
rect 2350 1118 11505 1137
rect 2794 1116 11505 1118
rect 9246 858 9349 873
rect 5511 842 5567 845
rect 2253 832 5567 842
rect 2253 798 5522 832
rect 5556 798 5567 832
rect 2253 788 5567 798
rect 9246 806 9271 858
rect 9323 806 9349 858
rect 9246 790 9349 806
rect 5511 786 5567 788
rect 497 679 560 685
rect 497 627 501 679
rect 553 627 560 679
rect 2369 667 2430 674
rect 2794 667 11510 668
rect 2369 634 11510 667
rect 2369 525 2979 634
rect 2373 518 2979 525
rect 3223 624 11510 634
rect 3223 572 11409 624
rect 11461 572 11510 624
rect 3223 554 11510 572
rect 3223 518 9871 554
rect 2373 502 9871 518
rect 9923 502 11510 554
rect 2373 499 11510 502
rect 2794 489 11510 499
rect 2811 316 2862 332
rect 2811 306 2818 316
rect 2782 286 2818 306
rect 2782 234 2795 286
rect 2852 282 2862 316
rect 2847 234 2862 282
rect 5108 322 5430 338
rect 5108 288 5114 322
rect 5148 288 5430 322
rect 7972 322 8172 338
rect 7972 320 8126 322
rect 5108 278 5430 288
rect 6741 310 6868 317
rect 6741 305 6803 310
rect 5108 272 5164 278
rect 6741 253 6779 305
rect 6837 276 6868 310
rect 6831 253 6868 276
rect 7962 316 8126 320
rect 7962 282 7978 316
rect 8012 288 8126 316
rect 8160 288 8172 322
rect 8012 282 8172 288
rect 7962 276 8172 282
rect 7962 268 8008 276
rect 8110 272 8172 276
rect 10413 316 10517 338
rect 10413 282 10423 316
rect 10457 313 10517 316
rect 6741 240 6868 253
rect 10413 261 10441 282
rect 10493 261 10517 313
rect 10413 238 10517 261
rect 2782 214 2862 234
rect 10454 41 10573 42
rect 2794 19 10573 41
rect 2794 -5 8278 19
rect 2794 -55 3770 -5
rect 3697 -185 3770 -55
rect 4078 -33 8278 -5
rect 8330 -33 8342 19
rect 8394 -33 8406 19
rect 8458 -33 8470 19
rect 8522 -33 8534 19
rect 8586 -33 8598 19
rect 8650 17 10573 19
rect 8650 -33 9552 17
rect 4078 -35 9552 -33
rect 9604 -35 9616 17
rect 9668 -35 10573 17
rect 4078 -55 10573 -35
rect 4078 -185 4153 -55
rect 10454 -56 10573 -55
rect 10419 -137 10795 -104
rect 3697 -251 4153 -185
rect 4321 -162 10795 -137
rect 4321 -163 10488 -162
rect 4321 -215 4461 -163
rect 4513 -215 10488 -163
rect 4321 -275 10488 -215
rect 4334 -578 4472 -275
rect 10419 -278 10488 -275
rect 10732 -278 10795 -162
rect 10419 -338 10795 -278
rect 16301 -122 16490 -104
rect 16301 -366 16337 -122
rect 16453 -366 16490 -122
rect 16301 -388 16490 -366
rect 3538 -716 4472 -578
rect 17158 -622 17417 -621
rect 9843 -663 9965 -653
rect 9843 -715 9846 -663
rect 9898 -715 9910 -663
rect 9962 -715 9965 -663
rect 17158 -674 17165 -622
rect 17217 -674 17229 -622
rect 17281 -674 17293 -622
rect 17345 -674 17357 -622
rect 17409 -674 17417 -622
rect 3538 -870 3676 -716
rect 9843 -724 9965 -715
rect 2647 -1008 3676 -870
rect 4464 -1014 6328 -833
rect 6147 -1316 6328 -1014
rect 16780 -1169 16928 -1164
rect 9553 -1207 9670 -1198
rect 9605 -1259 9617 -1207
rect 9669 -1259 9670 -1207
rect 16780 -1221 16796 -1169
rect 16848 -1221 16860 -1169
rect 16912 -1221 16928 -1169
rect 16780 -1225 16928 -1221
rect 9553 -1267 9670 -1259
rect 6147 -1356 7818 -1316
rect 6147 -1472 7596 -1356
rect 7776 -1472 7818 -1356
rect 6147 -1497 7818 -1472
rect 7529 -1508 7818 -1497
<< via1 >>
rect 2643 1366 2695 1375
rect 2643 1332 2653 1366
rect 2653 1332 2687 1366
rect 2687 1332 2695 1366
rect 2643 1323 2695 1332
rect 8279 1137 8331 1189
rect 8343 1137 8395 1189
rect 8407 1137 8459 1189
rect 8471 1137 8523 1189
rect 8535 1137 8587 1189
rect 8599 1137 8651 1189
rect 10869 1139 10921 1191
rect 10933 1139 10985 1191
rect 10997 1139 11049 1191
rect 9271 854 9323 858
rect 9271 820 9276 854
rect 9276 820 9310 854
rect 9310 820 9323 854
rect 9271 806 9323 820
rect 501 627 553 679
rect 2979 518 3223 634
rect 11409 572 11461 624
rect 9871 502 9923 554
rect 2795 282 2818 286
rect 2818 282 2847 286
rect 2795 234 2847 282
rect 6779 276 6803 305
rect 6803 276 6831 305
rect 6779 253 6831 276
rect 10441 282 10457 313
rect 10457 282 10493 313
rect 10441 261 10493 282
rect 3770 -185 4078 -5
rect 8278 -33 8330 19
rect 8342 -33 8394 19
rect 8406 -33 8458 19
rect 8470 -33 8522 19
rect 8534 -33 8586 19
rect 8598 -33 8650 19
rect 9552 -35 9604 17
rect 9616 -35 9668 17
rect 4461 -215 4513 -163
rect 10488 -278 10732 -162
rect 16337 -366 16453 -122
rect 9846 -715 9898 -663
rect 9910 -715 9962 -663
rect 17165 -674 17217 -622
rect 17229 -674 17281 -622
rect 17293 -674 17345 -622
rect 17357 -674 17409 -622
rect 9553 -1259 9605 -1207
rect 9617 -1259 9669 -1207
rect 16796 -1221 16848 -1169
rect 16860 -1221 16912 -1169
rect 7596 -1472 7776 -1356
<< metal2 >>
rect -7972 7723 25640 7992
rect -7972 5987 23832 7723
rect 25328 5987 25640 7723
rect -7972 5584 25640 5987
rect -6490 4978 22980 5277
rect -6490 3722 21607 4978
rect 22623 3722 22980 4978
rect -6490 3450 22980 3722
rect 10858 1804 12051 1981
rect 1817 1375 7256 1395
rect 1817 1323 2643 1375
rect 2695 1323 7256 1375
rect 1817 1308 7256 1323
rect 2611 1303 2727 1308
rect -973 832 -6 836
rect -973 789 4 832
rect -973 722 882 789
rect -973 648 4 722
rect -9109 278 4 648
rect -15673 -698 -15296 -697
rect -9109 -698 -8739 278
rect -973 275 4 278
rect 197 681 334 684
rect 496 681 562 685
rect 197 679 563 681
rect 197 627 501 679
rect 553 627 563 679
rect 197 622 563 627
rect -15673 -1068 -8739 -698
rect -15673 -1935 -15296 -1068
rect 197 -1438 334 622
rect 815 592 882 722
rect 1501 630 1874 697
rect 2934 644 3270 668
rect 2934 634 2993 644
rect 3209 634 3270 644
rect 1501 592 1568 630
rect 815 525 1568 592
rect 2934 518 2979 634
rect 3223 518 3270 634
rect 2934 508 2993 518
rect 3209 508 3270 518
rect 2934 488 3270 508
rect 4441 306 4539 308
rect 2782 286 4539 306
rect 2782 234 2795 286
rect 2847 234 4539 286
rect 6741 305 6868 317
rect 6741 253 6779 305
rect 6831 253 6868 305
rect 6741 240 6868 253
rect 2782 208 4539 234
rect 3697 -5 4153 39
rect 3697 -185 3770 -5
rect 4078 -185 4153 -5
rect 3697 -251 4153 -185
rect 4441 -163 4539 208
rect 6825 230 6868 240
rect 7191 230 7234 1308
rect 6825 187 7234 230
rect 8246 1189 8682 1212
rect 8246 1137 8279 1189
rect 8331 1137 8343 1189
rect 8395 1137 8407 1189
rect 8459 1137 8471 1189
rect 8523 1137 8535 1189
rect 8587 1137 8599 1189
rect 8651 1137 8682 1189
rect 8246 19 8682 1137
rect 10858 1191 11065 1804
rect 12384 1751 12524 1774
rect 12384 1695 12386 1751
rect 12442 1695 12466 1751
rect 12522 1695 12524 1751
rect 12384 1672 12524 1695
rect 17147 1710 17446 1784
rect 17147 1654 17176 1710
rect 17232 1654 17256 1710
rect 17312 1654 17336 1710
rect 17392 1654 17446 1710
rect 12410 1386 12713 1434
rect 12410 1250 12455 1386
rect 12671 1250 12713 1386
rect 12410 1199 12713 1250
rect 10858 1139 10869 1191
rect 10921 1139 10933 1191
rect 10985 1139 10997 1191
rect 11049 1139 11065 1191
rect 10858 1116 11065 1139
rect 9202 875 9352 919
rect 9202 819 9247 875
rect 9303 858 9352 875
rect 9202 806 9271 819
rect 9323 806 9352 858
rect 9202 775 9352 806
rect 11900 680 12051 720
rect 12780 719 16945 1207
rect 11369 624 11817 669
rect 9831 554 9975 578
rect 9831 502 9871 554
rect 9923 502 9975 554
rect 11369 572 11409 624
rect 11461 572 11817 624
rect 11900 624 11907 680
rect 11963 624 11987 680
rect 12043 624 12051 680
rect 11900 585 12051 624
rect 11369 523 11817 572
rect 8246 -33 8278 19
rect 8330 -33 8342 19
rect 8394 -33 8406 19
rect 8458 -33 8470 19
rect 8522 -33 8534 19
rect 8586 -33 8598 19
rect 8650 -33 8682 19
rect 8246 -55 8682 -33
rect 9542 17 9686 38
rect 9542 -35 9552 17
rect 9604 -35 9616 17
rect 9668 -35 9686 17
rect 4441 -215 4461 -163
rect 4513 -215 4539 -163
rect 4441 -241 4539 -215
rect 7759 -984 8238 -941
rect 4391 -1059 4723 -1036
rect 4391 -1195 4407 -1059
rect 4703 -1195 4723 -1059
rect 4391 -1219 4723 -1195
rect 7759 -1200 7819 -984
rect 8195 -1200 8238 -984
rect 7759 -1243 8238 -1200
rect 9542 -1207 9686 -35
rect 9831 -663 9975 502
rect 10417 315 10517 338
rect 10417 259 10439 315
rect 10495 259 10517 315
rect 10417 238 10517 259
rect 10987 134 11192 157
rect 10987 -2 11023 134
rect 11159 -2 11192 134
rect 15876 140 16098 174
rect 10987 -28 11192 -2
rect 11535 -25 12347 5
rect 15876 4 15920 140
rect 16056 4 16098 140
rect 15876 -22 16098 4
rect 11535 -81 11582 -25
rect 11638 -26 12347 -25
rect 11638 -81 12193 -26
rect 11535 -82 12193 -81
rect 12249 -82 12273 -26
rect 12329 -82 12347 -26
rect 10419 -152 10795 -104
rect 11535 -115 12347 -82
rect 10419 -288 10462 -152
rect 10758 -288 10795 -152
rect 10419 -338 10795 -288
rect 16301 -122 16490 -104
rect 16301 -136 16337 -122
rect 16453 -136 16490 -122
rect 16301 -352 16327 -136
rect 16463 -352 16490 -136
rect 16301 -366 16337 -352
rect 16453 -366 16490 -352
rect 16301 -388 16490 -366
rect 9831 -715 9846 -663
rect 9898 -715 9910 -663
rect 9962 -715 9975 -663
rect 9831 -740 9975 -715
rect 11806 -689 11842 -633
rect 11898 -689 11934 -633
rect 11806 -713 11934 -689
rect 11806 -769 11842 -713
rect 11898 -769 11934 -713
rect 15128 -794 15549 -740
rect 14913 -952 15098 -825
rect 15128 -1090 15197 -794
rect 15493 -1090 15549 -794
rect 15128 -1143 15549 -1090
rect 9542 -1259 9553 -1207
rect 9605 -1259 9617 -1207
rect 9669 -1259 9686 -1207
rect 16763 -1169 16945 719
rect 17147 -622 17446 1654
rect 18482 -475 18580 -436
rect 18482 -531 18503 -475
rect 18559 -531 18580 -475
rect 18482 -570 18580 -531
rect 17147 -674 17165 -622
rect 17217 -674 17229 -622
rect 17281 -674 17293 -622
rect 17345 -674 17357 -622
rect 17409 -674 17446 -622
rect 17147 -691 17446 -674
rect 16763 -1221 16796 -1169
rect 16848 -1221 16860 -1169
rect 16912 -1221 16945 -1169
rect 16763 -1246 16945 -1221
rect 9542 -1280 9686 -1259
rect 7555 -1346 7818 -1316
rect 7555 -1356 7618 -1346
rect 7754 -1356 7818 -1346
rect 247 -1439 302 -1438
rect 7555 -1472 7596 -1356
rect 7776 -1472 7818 -1356
rect 9226 -1357 9352 -1332
rect 9226 -1413 9261 -1357
rect 9317 -1413 9352 -1357
rect 9226 -1437 9352 -1413
rect 17747 -1359 17866 -1337
rect 17747 -1415 17778 -1359
rect 17834 -1415 17866 -1359
rect 17747 -1436 17866 -1415
rect 7555 -1482 7618 -1472
rect 7754 -1482 7818 -1472
rect 7555 -1508 7818 -1482
rect -6553 -8957 22930 -8773
rect -6553 -10453 21467 -8957
rect 22803 -10453 22930 -8957
rect -6553 -10600 22930 -10453
rect -7884 -11317 25640 -11076
rect -7884 -13133 23827 -11317
rect 25403 -13133 25640 -11317
rect -7884 -13484 25640 -13133
<< via2 >>
rect 23832 5987 25328 7723
rect 21607 3722 22623 4978
rect 2993 634 3209 644
rect 2993 518 3209 634
rect 2993 508 3209 518
rect 3776 -163 4072 -27
rect 12386 1695 12442 1751
rect 12466 1695 12522 1751
rect 17176 1654 17232 1710
rect 17256 1654 17312 1710
rect 17336 1654 17392 1710
rect 12455 1250 12671 1386
rect 9247 858 9303 875
rect 9247 819 9271 858
rect 9271 819 9303 858
rect 11907 624 11963 680
rect 11987 624 12043 680
rect 4407 -1195 4703 -1059
rect 7819 -1200 8195 -984
rect 10439 313 10495 315
rect 10439 261 10441 313
rect 10441 261 10493 313
rect 10493 261 10495 313
rect 10439 259 10495 261
rect 11023 -2 11159 134
rect 15920 4 16056 140
rect 11582 -81 11638 -25
rect 12193 -82 12249 -26
rect 12273 -82 12329 -26
rect 10462 -162 10758 -152
rect 10462 -278 10488 -162
rect 10488 -278 10732 -162
rect 10732 -278 10758 -162
rect 10462 -288 10758 -278
rect 16327 -352 16337 -136
rect 16337 -352 16453 -136
rect 16453 -352 16463 -136
rect 11842 -689 11898 -633
rect 11842 -769 11898 -713
rect 15197 -1090 15493 -794
rect 18503 -531 18559 -475
rect 7618 -1356 7754 -1346
rect 7618 -1472 7754 -1356
rect 9261 -1413 9317 -1357
rect 17778 -1415 17834 -1359
rect 7618 -1482 7754 -1472
rect 21467 -10453 22803 -8957
rect 23827 -13133 25403 -11317
<< metal3 >>
rect 23590 7723 25620 8020
rect 23590 5987 23832 7723
rect 25328 5987 25620 7723
rect 21330 4978 22950 5270
rect 21330 3722 21607 4978
rect 22623 3722 22950 4978
rect 12377 1751 17449 1784
rect 12377 1695 12386 1751
rect 12442 1695 12466 1751
rect 12522 1710 17449 1751
rect 12522 1695 17176 1710
rect 12377 1654 17176 1695
rect 17232 1654 17256 1710
rect 17312 1654 17336 1710
rect 17392 1654 17449 1710
rect 12377 1574 17449 1654
rect 12410 1386 12713 1434
rect 12410 1250 12455 1386
rect 12671 1309 12713 1386
rect 12671 1250 17672 1309
rect 12410 1137 17672 1250
rect 9202 875 9352 919
rect 9202 819 9247 875
rect 9303 819 9352 875
rect 9202 775 9352 819
rect 11791 735 11977 736
rect 11791 731 12059 735
rect 11791 680 12060 731
rect 2934 644 3270 665
rect 2934 508 2993 644
rect 3209 508 3270 644
rect 2934 -713 3270 508
rect 11791 624 11907 680
rect 11963 624 11987 680
rect 12043 624 12060 680
rect 11791 588 12060 624
rect 11791 572 12059 588
rect 10145 315 10517 338
rect 10145 259 10439 315
rect 10495 259 10517 315
rect 10145 238 10517 259
rect 3697 -23 4153 39
rect 3697 -167 3772 -23
rect 4076 -167 4153 -23
rect 3697 -251 4153 -167
rect 10145 -445 10245 238
rect 10990 138 11191 157
rect 10990 -6 11019 138
rect 11163 -6 11191 138
rect 10990 -22 11191 -6
rect 11535 -25 11685 4
rect 11535 -81 11582 -25
rect 11638 -81 11685 -25
rect 11535 -104 11685 -81
rect 10419 -152 11687 -104
rect 10419 -288 10462 -152
rect 10758 -288 11687 -152
rect 10419 -338 11687 -288
rect 10145 -545 11518 -445
rect 7759 -984 8238 -941
rect 4391 -1055 4723 -1036
rect 4391 -1059 4443 -1055
rect 4667 -1059 4723 -1055
rect 4391 -1195 4407 -1059
rect 4703 -1195 4723 -1059
rect 4391 -1199 4443 -1195
rect 4667 -1199 4723 -1195
rect 4391 -1219 4723 -1199
rect 7759 -1200 7819 -984
rect 8195 -1200 8238 -984
rect 7759 -1243 8238 -1200
rect 7555 -1342 7818 -1316
rect 11418 -1319 11518 -545
rect 11791 -633 11977 572
rect 15876 144 16098 174
rect 12177 -26 12348 23
rect 15876 0 15916 144
rect 16060 0 16098 144
rect 15876 -22 16098 0
rect 12177 -82 12193 -26
rect 12249 -82 12273 -26
rect 12329 -82 12348 -26
rect 12177 -104 12348 -82
rect 12177 -127 16490 -104
rect 12180 -136 16490 -127
rect 12180 -338 16327 -136
rect 16301 -352 16327 -338
rect 16463 -352 16490 -136
rect 16301 -388 16490 -352
rect 17500 -267 17672 1137
rect 17500 -416 18381 -267
rect 17500 -439 18598 -416
rect 18209 -475 18598 -439
rect 18209 -531 18503 -475
rect 18559 -531 18598 -475
rect 18209 -588 18598 -531
rect 11791 -689 11842 -633
rect 11898 -689 11977 -633
rect 11791 -713 11977 -689
rect 11791 -769 11842 -713
rect 11898 -769 11977 -713
rect 11791 -787 11977 -769
rect 11791 -788 11950 -787
rect 15128 -790 15549 -740
rect 15128 -1094 15193 -790
rect 15497 -1094 15549 -790
rect 15128 -1143 15549 -1094
rect 7555 -1486 7614 -1342
rect 7758 -1486 7818 -1342
rect 9216 -1352 17879 -1319
rect 9216 -1416 9253 -1352
rect 9317 -1359 17879 -1352
rect 9317 -1415 17778 -1359
rect 17834 -1415 17879 -1359
rect 9317 -1416 17879 -1415
rect 9216 -1452 17879 -1416
rect 7555 -1508 7818 -1486
rect 6877 -1875 7364 -1669
rect 6877 -2059 7083 -1875
rect 5254 -2265 7085 -2059
rect 21330 -8957 22950 3722
rect 21330 -10453 21467 -8957
rect 22803 -10453 22950 -8957
rect 21330 -10600 22950 -10453
rect 23590 -11317 25620 5987
rect 23590 -13133 23827 -11317
rect 25403 -13133 25620 -11317
rect 23590 -13400 25620 -13133
<< via3 >>
rect 3772 -27 4076 -23
rect 3772 -163 3776 -27
rect 3776 -163 4072 -27
rect 4072 -163 4076 -27
rect 3772 -167 4076 -163
rect 11019 134 11163 138
rect 11019 -2 11023 134
rect 11023 -2 11159 134
rect 11159 -2 11163 134
rect 11019 -6 11163 -2
rect 4443 -1059 4667 -1055
rect 4443 -1195 4667 -1059
rect 4443 -1199 4667 -1195
rect 15916 140 16060 144
rect 15916 4 15920 140
rect 15920 4 16056 140
rect 16056 4 16060 140
rect 15916 0 16060 4
rect 15193 -794 15497 -790
rect 15193 -1090 15197 -794
rect 15197 -1090 15493 -794
rect 15493 -1090 15497 -794
rect 15193 -1094 15497 -1090
rect 7614 -1346 7758 -1342
rect 7614 -1482 7618 -1346
rect 7618 -1482 7754 -1346
rect 7754 -1482 7758 -1346
rect 7614 -1486 7758 -1482
rect 9253 -1357 9317 -1352
rect 9253 -1413 9261 -1357
rect 9261 -1413 9317 -1357
rect 9253 -1416 9317 -1413
<< metal4 >>
rect 10990 155 11191 157
rect 15876 155 16098 174
rect 10990 144 16098 155
rect 10990 138 15916 144
rect 3697 -23 4153 39
rect 10990 -6 11019 138
rect 11163 0 15916 138
rect 16060 0 16098 144
rect 11163 -6 16098 0
rect 10990 -22 16098 -6
rect 10990 -23 16097 -22
rect 3697 -167 3772 -23
rect 4076 -167 4153 -23
rect 3697 -251 4153 -167
rect 11440 -383 11618 -23
rect 5327 -561 11618 -383
rect 5327 -1035 5505 -561
rect 4391 -1055 5505 -1035
rect 4391 -1199 4443 -1055
rect 4667 -1199 5505 -1055
rect 15128 -790 15549 -740
rect 15128 -1094 15193 -790
rect 15497 -1094 15549 -790
rect 15128 -1143 15549 -1094
rect 4391 -1213 5505 -1199
rect 4391 -1219 4723 -1213
rect 7555 -1342 9366 -1316
rect 7555 -1486 7614 -1342
rect 7758 -1352 9366 -1342
rect 7758 -1416 9253 -1352
rect 9317 -1416 9366 -1352
rect 7758 -1486 9366 -1416
rect 7555 -1506 9366 -1486
rect 7555 -1508 7818 -1506
rect -5611 -5077 -3460 -4669
rect -5611 -6913 -5306 -5077
rect -3790 -6913 -3460 -5077
rect -5611 -7399 -3460 -6913
<< via4 >>
rect 15227 -1060 15463 -824
rect -5306 -6913 -3790 -5077
<< metal5 >>
rect 15127 -824 15549 -740
rect 15127 -1060 15227 -824
rect 15463 -1060 15549 -824
rect 15127 -1143 15549 -1060
rect -5611 -4684 -3460 -4669
rect 15127 -4684 15539 -1143
rect -5611 -5077 15539 -4684
rect -5611 -6913 -5306 -5077
rect -3790 -5140 15539 -5077
rect -3790 -6913 -3460 -5140
rect -5611 -7399 -3460 -6913
use COMPA  COMPA_0
timestamp 1667803582
transform -1 0 2295 0 1 100
box -186 -194 2295 1896
use DAC  DAC_0
timestamp 1667803582
transform 1 0 11854 0 1 879
box -2619 -720 977 1200
use Delay_Block  Delay_Block_0
timestamp 1667803582
transform 1 0 2794 0 1 620
box -38 -48 2447 592
use Integrator_n  Integrator_n_0
timestamp 1667803582
transform -1 0 -391 0 1 -13484
box -6976 0 30217 21478
use NOCFINAL  NOCFINAL_0
timestamp 1667803582
transform -1 0 6807 0 -1 535
box -1270 -50 1608 592
use Subtractor_Mag  Subtractor_Mag_0
timestamp 1667803582
transform 1 0 15836 0 1 -2197
box -1952 -5933 4099 2586
use Subtractor_Mag  Subtractor_Mag_1
timestamp 1667803582
transform -1 0 11260 0 1 -2235
box -1952 -5933 4099 2586
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_0
timestamp 1667803582
transform 1 0 6743 0 1 620
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_1
timestamp 1667803582
transform 1 0 8089 0 -1 537
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_2
timestamp 1667803582
transform -1 0 5186 0 -1 537
box -38 -48 2430 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0
timestamp 1667803582
transform 1 0 5237 0 1 620
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1667803582
transform -1 0 10573 0 -1 537
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1667803582
transform 1 0 9135 0 1 620
box -38 -48 130 592
<< labels >>
flabel metal2 s 8377 1179 8377 1179 0 FreeSans 4000 0 0 0 VDD
port 1 nsew
flabel metal1 s 9826 576 9826 576 0 FreeSans 4000 0 0 0 VSS
port 2 nsew
flabel metal3 s 7987 -1069 7987 -1069 0 FreeSans 3000 0 0 0 SD_IN_1
port 3 nsew
flabel metal2 s 3234 1363 3234 1363 0 FreeSans 8000 0 0 0 CLK
port 4 nsew
flabel metal3 s 9259 863 9259 863 0 FreeSans 3000 0 0 0 SD_DOUT_1
port 5 nsew
<< end >>
