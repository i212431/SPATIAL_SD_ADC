magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< nwell >>
rect 433 1466 1546 1758
rect -53 728 2019 1466
<< metal1 >>
rect -134 1798 2056 1874
rect -134 994 -58 1798
rect 226 1748 2056 1798
rect -12 960 131 1736
rect 185 1725 2056 1748
rect 185 1688 2059 1725
rect 185 1421 446 1688
rect 498 1598 610 1599
rect 498 1422 762 1598
rect 185 1407 443 1421
rect 538 1410 542 1422
rect 185 1397 432 1407
rect 349 1076 393 1397
rect 440 1274 507 1369
rect 440 1222 444 1274
rect 496 1222 507 1274
rect 440 1116 507 1222
rect 598 1166 634 1422
rect 816 1421 851 1688
rect 908 1496 1006 1524
rect 908 1444 929 1496
rect 981 1444 1006 1496
rect 908 1410 1006 1444
rect 1389 1420 1422 1688
rect 1475 1489 1743 1595
rect 1475 1437 1507 1489
rect 1559 1437 1743 1489
rect 1475 1423 1743 1437
rect 910 1369 990 1410
rect 1478 1408 1626 1423
rect 1795 1416 2056 1688
rect 757 1298 990 1369
rect 570 1132 662 1166
rect 570 1080 592 1132
rect 644 1080 662 1132
rect -125 23 -78 537
rect -12 481 42 960
rect 113 886 223 915
rect 113 834 141 886
rect 193 834 223 886
rect 349 872 452 1076
rect 502 840 537 1062
rect 541 888 542 1076
rect 570 1052 662 1080
rect 757 1059 935 1298
rect 1300 1135 1485 1368
rect 1300 1083 1340 1135
rect 1392 1083 1485 1135
rect 598 971 634 1052
rect 757 1008 936 1059
rect 593 954 675 971
rect 593 902 616 954
rect 668 902 675 954
rect 593 891 675 902
rect 598 888 675 891
rect 113 808 223 834
rect 124 527 191 808
rect 501 799 577 840
rect 501 723 647 799
rect 417 591 525 603
rect 417 539 446 591
rect 498 539 525 591
rect 417 527 525 539
rect 571 486 647 723
rect 758 688 936 1008
rect 1300 1006 1485 1083
rect 764 529 936 688
rect 964 932 1040 978
rect 964 880 971 932
rect 1023 880 1040 932
rect 1303 957 1367 1006
rect 1549 963 1626 1408
rect 1734 1274 1801 1371
rect 1734 1222 1740 1274
rect 1792 1222 1801 1274
rect 1734 1119 1801 1222
rect 1891 1063 1946 1416
rect 1303 893 1415 957
rect 964 844 1040 880
rect 964 496 1013 844
rect 1210 779 1279 792
rect 1210 727 1218 779
rect 1270 727 1279 779
rect 1210 719 1279 727
rect -12 106 131 481
rect -12 105 42 106
rect 184 23 231 483
rect 571 448 867 486
rect 501 407 867 448
rect 925 411 1013 496
rect 1079 686 1164 698
rect 1079 634 1095 686
rect 1147 634 1164 686
rect 501 377 650 407
rect 571 372 647 377
rect 383 198 448 254
rect 383 146 392 198
rect 444 146 448 198
rect 1079 173 1164 634
rect 1213 497 1252 719
rect 1351 592 1415 893
rect 1478 947 1626 963
rect 1478 895 1484 947
rect 1536 895 1626 947
rect 1478 883 1626 895
rect 1699 827 1744 1063
rect 1795 886 1946 1063
rect 2104 953 2267 1733
rect 2050 859 2113 906
rect 1307 528 1415 592
rect 1615 768 1746 827
rect 2050 807 2058 859
rect 2110 807 2113 859
rect 1615 519 1674 768
rect 1733 526 1806 575
rect 2050 527 2113 807
rect 1212 408 1304 497
rect 1615 483 1702 519
rect 2189 483 2267 953
rect 1362 480 1702 483
rect 1362 377 1744 480
rect 1615 322 1744 377
rect 1243 184 1335 213
rect 383 104 448 146
rect 1243 132 1260 184
rect 1312 132 1335 184
rect 1243 44 1335 132
rect 1795 197 1869 238
rect 1795 145 1801 197
rect 1853 145 1869 197
rect 1795 104 1869 145
rect -125 -91 1076 23
rect 1129 -48 1335 44
rect 2011 23 2056 481
rect 2104 103 2267 483
rect 1402 -91 2056 23
rect -125 -100 2056 -91
rect 1038 -125 1454 -100
<< via1 >>
rect 444 1222 496 1274
rect 929 1444 981 1496
rect 1507 1437 1559 1489
rect 592 1080 644 1132
rect 141 834 193 886
rect 1340 1083 1392 1135
rect 616 902 668 954
rect 446 539 498 591
rect 971 880 1023 932
rect 1740 1222 1792 1274
rect 1218 727 1270 779
rect 1095 634 1147 686
rect 392 146 444 198
rect 1484 895 1536 947
rect 2058 807 2110 859
rect 1260 132 1312 184
rect 1801 145 1853 197
<< metal2 >>
rect 910 1496 1584 1522
rect 910 1444 929 1496
rect 981 1489 1584 1496
rect 981 1444 1507 1489
rect 910 1437 1507 1444
rect 1559 1437 1584 1489
rect 910 1408 1584 1437
rect 1077 1288 1164 1289
rect 436 1274 1801 1288
rect 436 1222 444 1274
rect 496 1222 1740 1274
rect 1792 1222 1801 1274
rect 436 1210 1801 1222
rect 570 1134 662 1166
rect 570 1078 590 1134
rect 646 1078 662 1134
rect 570 1052 662 1078
rect 964 968 1040 978
rect 654 967 1040 968
rect 113 954 1040 967
rect 113 902 616 954
rect 668 932 1040 954
rect 668 902 971 932
rect 113 886 971 902
rect 113 834 141 886
rect 193 880 971 886
rect 1023 880 1040 932
rect 193 844 1040 880
rect 193 843 1012 844
rect 193 834 223 843
rect 113 808 223 834
rect 1077 686 1164 1210
rect 1302 1137 1428 1162
rect 1302 1081 1338 1137
rect 1394 1081 1428 1137
rect 1302 1064 1428 1081
rect 1471 947 2115 959
rect 1471 895 1484 947
rect 1536 895 2115 947
rect 1471 890 2115 895
rect 1212 859 2115 890
rect 1212 807 2058 859
rect 2110 807 2115 859
rect 1212 799 2115 807
rect 1212 792 1303 799
rect 1210 779 1303 792
rect 1210 727 1218 779
rect 1270 727 1303 779
rect 1210 723 1303 727
rect 1210 719 1279 723
rect 1077 634 1095 686
rect 1147 634 1164 686
rect 1077 622 1164 634
rect 417 591 525 603
rect 417 539 446 591
rect 498 539 525 591
rect 417 527 525 539
rect 1248 236 1355 237
rect 382 198 1870 236
rect 382 146 392 198
rect 444 197 1870 198
rect 444 184 1801 197
rect 444 146 1260 184
rect 382 132 1260 146
rect 1312 145 1801 184
rect 1853 145 1870 197
rect 1312 132 1870 145
rect 382 104 1870 132
<< via2 >>
rect 590 1132 646 1134
rect 590 1080 592 1132
rect 592 1080 644 1132
rect 644 1080 646 1132
rect 590 1078 646 1080
rect 1338 1135 1394 1137
rect 1338 1083 1340 1135
rect 1340 1083 1392 1135
rect 1392 1083 1394 1135
rect 1338 1081 1394 1083
<< metal3 >>
rect 570 1162 662 1166
rect 570 1137 1426 1162
rect 570 1134 1338 1137
rect 570 1078 590 1134
rect 646 1081 1338 1134
rect 1394 1081 1426 1137
rect 646 1078 1426 1081
rect 570 1062 1426 1078
rect 570 1052 662 1062
use sky130_fd_pr__nfet_01v8_6H5H3D  sky130_fd_pr__nfet_01v8_6H5H3D_0
timestamp 1667803582
transform 1 0 2079 0 1 327
box -201 -369 201 369
use sky130_fd_pr__nfet_01v8_6H5H3D  sky130_fd_pr__nfet_01v8_6H5H3D_1
timestamp 1667803582
transform 1 0 1768 0 1 327
box -201 -369 201 369
use sky130_fd_pr__nfet_01v8_6H5H3D  sky130_fd_pr__nfet_01v8_6H5H3D_2
timestamp 1667803582
transform 1 0 474 0 1 326
box -201 -369 201 369
use sky130_fd_pr__nfet_01v8_6H5H3D  sky130_fd_pr__nfet_01v8_6H5H3D_3
timestamp 1667803582
transform 1 0 158 0 1 326
box -201 -369 201 369
use sky130_fd_pr__nfet_01v8_LDKBCP  sky130_fd_pr__nfet_01v8_LDKBCP_0
timestamp 1667803582
transform 1 0 1335 0 1 476
box -201 -219 201 219
use sky130_fd_pr__nfet_01v8_LDKBCP  sky130_fd_pr__nfet_01v8_LDKBCP_1
timestamp 1667803582
transform 1 0 896 0 1 477
box -201 -219 201 219
use sky130_fd_pr__nfet_01v8_RB5HKB  sky130_fd_pr__nfet_01v8_RB5HKB_0
timestamp 1667803582
transform 1 0 1103 0 1 75
box -201 -269 201 269
use sky130_fd_pr__pfet_01v8_LTABJ9  sky130_fd_pr__pfet_01v8_LTABJ9_0
timestamp 1667803582
transform 1 0 2084 0 1 1312
box -211 -584 211 584
use sky130_fd_pr__pfet_01v8_LTABJ9  sky130_fd_pr__pfet_01v8_LTABJ9_1
timestamp 1667803582
transform 1 0 158 0 1 1312
box -211 -584 211 584
use sky130_fd_pr__pfet_01v8_LZABJ9  sky130_fd_pr__pfet_01v8_LZABJ9_0
timestamp 1667803582
transform -1 0 1768 0 -1 1012
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_LZABJ9  sky130_fd_pr__pfet_01v8_LZABJ9_1
timestamp 1667803582
transform 1 0 1768 0 1 1474
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_LZABJ9  sky130_fd_pr__pfet_01v8_LZABJ9_2
timestamp 1667803582
transform 1 0 1452 0 1 1474
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_LZABJ9  sky130_fd_pr__pfet_01v8_LZABJ9_3
timestamp 1667803582
transform 1 0 474 0 1 1474
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_LZABJ9  sky130_fd_pr__pfet_01v8_LZABJ9_4
timestamp 1667803582
transform -1 0 474 0 -1 1012
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_LZABJ9  sky130_fd_pr__pfet_01v8_LZABJ9_5
timestamp 1667803582
transform 1 0 790 0 1 1474
box -211 -284 211 284
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1667803582
transform 1 0 -148 0 1 488
box -38 -48 130 592
<< labels >>
flabel metal1 s 15 709 15 709 0 FreeSans 800 0 0 0 VOUTP
port 1 nsew
flabel metal1 s 1050 1773 1050 1773 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal1 s 2233 711 2233 711 0 FreeSans 800 0 0 0 VOUTN
port 3 nsew
flabel metal1 s 1768 550 1768 550 0 FreeSans 800 0 0 0 VINN
port 4 nsew
flabel metal2 s 1108 1255 1108 1255 0 FreeSans 800 0 0 0 CLK
port 5 nsew
flabel metal2 s 475 565 475 565 0 FreeSans 800 0 0 0 VINP
port 6 nsew
flabel metal1 s 662 -84 662 -84 0 FreeSans 1200 0 0 0 VSS
port 7 nsew
<< end >>
