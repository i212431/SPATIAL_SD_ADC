magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< nwell >>
rect -50 1383 -20 1881
rect -50 1040 478 1383
rect -511 942 478 1040
rect -490 757 478 942
rect -227 719 14 757
<< poly >>
rect 62 1845 398 1916
rect 44 722 380 793
rect 62 609 398 676
rect 44 0 380 66
<< locali >>
rect -551 895 -517 909
rect -551 823 -517 861
rect -551 776 -517 789
<< viali >>
rect -551 861 -517 895
rect -551 789 -517 823
<< metal1 >>
rect 62 1860 541 1906
rect -8 1753 61 1781
rect -8 1701 0 1753
rect 52 1701 61 1753
rect -8 1689 61 1701
rect -8 1637 0 1689
rect 52 1637 61 1689
rect -8 1609 61 1637
rect 188 1752 254 1781
rect 188 1700 195 1752
rect 247 1700 254 1752
rect 188 1688 254 1700
rect 188 1636 195 1688
rect 247 1636 254 1688
rect 188 1609 254 1636
rect 380 1753 453 1781
rect 380 1701 390 1753
rect 442 1701 453 1753
rect 380 1689 453 1701
rect 380 1637 390 1689
rect 442 1637 453 1689
rect 380 1609 453 1637
rect 91 1051 158 1071
rect -2604 954 -248 1050
rect 91 999 98 1051
rect 150 999 158 1051
rect 91 987 158 999
rect 91 935 98 987
rect 150 935 158 987
rect 91 923 158 935
rect -560 895 -509 921
rect -560 861 -551 895
rect -517 861 -509 895
rect -560 823 -509 861
rect 91 871 98 923
rect 150 871 158 923
rect 91 851 158 871
rect 284 1051 351 1071
rect 284 999 291 1051
rect 343 999 351 1051
rect 284 987 351 999
rect 284 935 291 987
rect 343 935 351 987
rect 284 923 351 935
rect 284 871 291 923
rect 343 871 351 923
rect 284 851 351 871
rect -560 789 -551 823
rect -517 789 -509 823
rect -560 778 -509 789
rect 495 778 541 1860
rect -560 772 541 778
rect -559 732 541 772
rect -758 699 -597 719
rect -758 666 -123 699
rect -758 653 541 666
rect -169 620 541 653
rect 91 527 159 556
rect -2604 410 -248 506
rect 91 475 98 527
rect 150 475 159 527
rect 91 463 159 475
rect 91 411 98 463
rect 150 411 159 463
rect 91 383 159 411
rect 284 527 351 556
rect 284 475 292 527
rect 344 475 351 527
rect 284 463 351 475
rect 284 411 292 463
rect 344 411 351 463
rect 284 383 351 411
rect -5 267 62 304
rect -5 215 1 267
rect 53 215 62 267
rect -5 203 62 215
rect -5 151 1 203
rect 53 151 62 203
rect -5 115 62 151
rect 188 266 254 303
rect 188 214 195 266
rect 247 214 254 266
rect 188 202 254 214
rect 188 150 195 202
rect 247 150 254 202
rect 188 115 254 150
rect 380 266 442 302
rect 380 214 384 266
rect 436 214 442 266
rect 380 202 442 214
rect 380 150 384 202
rect 436 150 442 202
rect 380 115 442 150
rect 495 56 541 620
rect 43 10 541 56
<< via1 >>
rect 0 1701 52 1753
rect 0 1637 52 1689
rect 195 1700 247 1752
rect 195 1636 247 1688
rect 390 1701 442 1753
rect 390 1637 442 1689
rect 98 999 150 1051
rect 98 935 150 987
rect 98 871 150 923
rect 291 999 343 1051
rect 291 935 343 987
rect 291 871 343 923
rect 98 475 150 527
rect 98 411 150 463
rect 292 475 344 527
rect 292 411 344 463
rect 1 215 53 267
rect 1 151 53 203
rect 195 214 247 266
rect 195 150 247 202
rect 384 214 436 266
rect 384 150 436 202
<< metal2 >>
rect -12 1753 453 1781
rect -12 1701 0 1753
rect 52 1752 390 1753
rect 52 1701 195 1752
rect -12 1700 195 1701
rect 247 1701 390 1752
rect 442 1701 453 1753
rect 247 1700 453 1701
rect -12 1689 453 1700
rect -12 1637 0 1689
rect 52 1688 390 1689
rect 52 1637 195 1688
rect -12 1636 195 1637
rect 247 1637 390 1688
rect 442 1637 453 1689
rect 247 1636 453 1637
rect -12 1609 453 1636
rect 91 1051 351 1071
rect 91 999 98 1051
rect 150 999 291 1051
rect 343 999 351 1051
rect 91 987 351 999
rect 91 935 98 987
rect 150 935 291 987
rect 343 935 351 987
rect 91 923 351 935
rect 91 871 98 923
rect 150 871 291 923
rect 343 871 351 923
rect 91 527 351 871
rect 91 475 98 527
rect 150 475 292 527
rect 344 475 351 527
rect 91 463 351 475
rect 91 411 98 463
rect 150 411 292 463
rect 344 411 351 463
rect 91 383 351 411
rect 380 303 442 1609
rect -5 267 442 303
rect -5 215 1 267
rect 53 266 442 267
rect 53 215 195 266
rect -5 214 195 215
rect 247 214 384 266
rect 436 214 442 266
rect -5 203 442 214
rect -5 151 1 203
rect 53 202 442 203
rect 53 151 195 202
rect -5 150 195 151
rect 247 150 384 202
rect 436 150 442 202
rect -5 115 442 150
use sky130_fd_pr__nfet_01v8_JRYMCH  sky130_fd_pr__nfet_01v8_JRYMCH_0
timestamp 1667803582
transform 1 0 221 0 1 338
box -247 -338 247 338
use sky130_fd_pr__pfet_01v8_52DJHB  sky130_fd_pr__pfet_01v8_52DJHB_0
timestamp 1667803582
transform 1 0 221 0 1 1319
box -257 -600 257 600
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0
timestamp 1667803582
transform 1 0 -2604 0 1 458
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1667803582
transform 1 0 -340 0 1 458
box -38 -48 130 592
<< labels >>
flabel metal2 s 419 698 419 698 0 FreeSans 1000 0 0 0 B
port 1 nsew
flabel metal2 s 177 704 177 704 0 FreeSans 1000 0 0 0 A
port 2 nsew
flabel metal1 s -538 823 -538 823 0 FreeSans 1000 0 0 0 CLKB
port 3 nsew
flabel metal1 s -1487 986 -1487 986 0 FreeSans 1000 0 0 0 VDD
port 4 nsew
flabel metal1 s -1466 440 -1466 440 0 FreeSans 1000 0 0 0 VSS
port 5 nsew
<< end >>
