magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< error_p >>
rect -29 -111 29 -105
rect -29 -145 -17 -111
rect -29 -151 29 -145
<< nwell >>
rect -211 -284 211 284
<< pmos >>
rect -15 -64 15 136
<< pdiff >>
rect -73 121 -15 136
rect -73 87 -61 121
rect -27 87 -15 121
rect -73 53 -15 87
rect -73 19 -61 53
rect -27 19 -15 53
rect -73 -15 -15 19
rect -73 -49 -61 -15
rect -27 -49 -15 -15
rect -73 -64 -15 -49
rect 15 121 73 136
rect 15 87 27 121
rect 61 87 73 121
rect 15 53 73 87
rect 15 19 27 53
rect 61 19 73 53
rect 15 -15 73 19
rect 15 -49 27 -15
rect 61 -49 73 -15
rect 15 -64 73 -49
<< pdiffc >>
rect -61 87 -27 121
rect -61 19 -27 53
rect -61 -49 -27 -15
rect 27 87 61 121
rect 27 19 61 53
rect 27 -49 61 -15
<< nsubdiff >>
rect -175 214 175 248
rect -175 -214 -141 214
rect 141 -214 175 214
rect -175 -248 175 -214
<< poly >>
rect -15 136 15 162
rect -15 -95 15 -64
rect -33 -111 33 -95
rect -33 -145 -17 -111
rect 17 -145 33 -111
rect -33 -161 33 -145
<< polycont >>
rect -17 -145 17 -111
<< locali >>
rect -175 214 175 248
rect -175 -214 -141 214
rect -61 121 -27 140
rect -61 53 -27 55
rect -61 17 -27 19
rect -61 -68 -27 -49
rect 27 121 61 140
rect 27 53 61 55
rect 27 17 61 19
rect 27 -68 61 -49
rect -33 -145 -17 -111
rect 17 -145 33 -111
rect 141 -214 175 214
rect -175 -248 175 -214
<< viali >>
rect -61 87 -27 89
rect -61 55 -27 87
rect -61 -15 -27 17
rect -61 -17 -27 -15
rect 27 87 61 89
rect 27 55 61 87
rect 27 -15 61 17
rect 27 -17 61 -15
rect -17 -145 17 -111
<< metal1 >>
rect -67 89 -21 136
rect -67 55 -61 89
rect -27 55 -21 89
rect -67 17 -21 55
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -64 -21 -17
rect 21 89 67 136
rect 21 55 27 89
rect 61 55 67 89
rect 21 17 67 55
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -64 67 -17
rect -29 -111 29 -105
rect -29 -145 -17 -111
rect 17 -145 29 -111
rect -29 -151 29 -145
<< properties >>
string FIXED_BBOX -158 -231 158 231
<< end >>
