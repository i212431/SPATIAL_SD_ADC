magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< metal3 >>
rect -2950 2872 2949 2900
rect -2950 2808 2865 2872
rect 2929 2808 2949 2872
rect -2950 2792 2949 2808
rect -2950 2728 2865 2792
rect 2929 2728 2949 2792
rect -2950 2712 2949 2728
rect -2950 2648 2865 2712
rect 2929 2648 2949 2712
rect -2950 2632 2949 2648
rect -2950 2568 2865 2632
rect 2929 2568 2949 2632
rect -2950 2552 2949 2568
rect -2950 2488 2865 2552
rect 2929 2488 2949 2552
rect -2950 2472 2949 2488
rect -2950 2408 2865 2472
rect 2929 2408 2949 2472
rect -2950 2392 2949 2408
rect -2950 2328 2865 2392
rect 2929 2328 2949 2392
rect -2950 2312 2949 2328
rect -2950 2248 2865 2312
rect 2929 2248 2949 2312
rect -2950 2232 2949 2248
rect -2950 2168 2865 2232
rect 2929 2168 2949 2232
rect -2950 2152 2949 2168
rect -2950 2088 2865 2152
rect 2929 2088 2949 2152
rect -2950 2072 2949 2088
rect -2950 2008 2865 2072
rect 2929 2008 2949 2072
rect -2950 1992 2949 2008
rect -2950 1928 2865 1992
rect 2929 1928 2949 1992
rect -2950 1912 2949 1928
rect -2950 1848 2865 1912
rect 2929 1848 2949 1912
rect -2950 1832 2949 1848
rect -2950 1768 2865 1832
rect 2929 1768 2949 1832
rect -2950 1752 2949 1768
rect -2950 1688 2865 1752
rect 2929 1688 2949 1752
rect -2950 1672 2949 1688
rect -2950 1608 2865 1672
rect 2929 1608 2949 1672
rect -2950 1592 2949 1608
rect -2950 1528 2865 1592
rect 2929 1528 2949 1592
rect -2950 1512 2949 1528
rect -2950 1448 2865 1512
rect 2929 1448 2949 1512
rect -2950 1432 2949 1448
rect -2950 1368 2865 1432
rect 2929 1368 2949 1432
rect -2950 1352 2949 1368
rect -2950 1288 2865 1352
rect 2929 1288 2949 1352
rect -2950 1272 2949 1288
rect -2950 1208 2865 1272
rect 2929 1208 2949 1272
rect -2950 1192 2949 1208
rect -2950 1128 2865 1192
rect 2929 1128 2949 1192
rect -2950 1112 2949 1128
rect -2950 1048 2865 1112
rect 2929 1048 2949 1112
rect -2950 1032 2949 1048
rect -2950 968 2865 1032
rect 2929 968 2949 1032
rect -2950 952 2949 968
rect -2950 888 2865 952
rect 2929 888 2949 952
rect -2950 872 2949 888
rect -2950 808 2865 872
rect 2929 808 2949 872
rect -2950 792 2949 808
rect -2950 728 2865 792
rect 2929 728 2949 792
rect -2950 712 2949 728
rect -2950 648 2865 712
rect 2929 648 2949 712
rect -2950 632 2949 648
rect -2950 568 2865 632
rect 2929 568 2949 632
rect -2950 552 2949 568
rect -2950 488 2865 552
rect 2929 488 2949 552
rect -2950 472 2949 488
rect -2950 408 2865 472
rect 2929 408 2949 472
rect -2950 392 2949 408
rect -2950 328 2865 392
rect 2929 328 2949 392
rect -2950 312 2949 328
rect -2950 248 2865 312
rect 2929 248 2949 312
rect -2950 232 2949 248
rect -2950 168 2865 232
rect 2929 168 2949 232
rect -2950 152 2949 168
rect -2950 88 2865 152
rect 2929 88 2949 152
rect -2950 72 2949 88
rect -2950 8 2865 72
rect 2929 8 2949 72
rect -2950 -8 2949 8
rect -2950 -72 2865 -8
rect 2929 -72 2949 -8
rect -2950 -88 2949 -72
rect -2950 -152 2865 -88
rect 2929 -152 2949 -88
rect -2950 -168 2949 -152
rect -2950 -232 2865 -168
rect 2929 -232 2949 -168
rect -2950 -248 2949 -232
rect -2950 -312 2865 -248
rect 2929 -312 2949 -248
rect -2950 -328 2949 -312
rect -2950 -392 2865 -328
rect 2929 -392 2949 -328
rect -2950 -408 2949 -392
rect -2950 -472 2865 -408
rect 2929 -472 2949 -408
rect -2950 -488 2949 -472
rect -2950 -552 2865 -488
rect 2929 -552 2949 -488
rect -2950 -568 2949 -552
rect -2950 -632 2865 -568
rect 2929 -632 2949 -568
rect -2950 -648 2949 -632
rect -2950 -712 2865 -648
rect 2929 -712 2949 -648
rect -2950 -728 2949 -712
rect -2950 -792 2865 -728
rect 2929 -792 2949 -728
rect -2950 -808 2949 -792
rect -2950 -872 2865 -808
rect 2929 -872 2949 -808
rect -2950 -888 2949 -872
rect -2950 -952 2865 -888
rect 2929 -952 2949 -888
rect -2950 -968 2949 -952
rect -2950 -1032 2865 -968
rect 2929 -1032 2949 -968
rect -2950 -1048 2949 -1032
rect -2950 -1112 2865 -1048
rect 2929 -1112 2949 -1048
rect -2950 -1128 2949 -1112
rect -2950 -1192 2865 -1128
rect 2929 -1192 2949 -1128
rect -2950 -1208 2949 -1192
rect -2950 -1272 2865 -1208
rect 2929 -1272 2949 -1208
rect -2950 -1288 2949 -1272
rect -2950 -1352 2865 -1288
rect 2929 -1352 2949 -1288
rect -2950 -1368 2949 -1352
rect -2950 -1432 2865 -1368
rect 2929 -1432 2949 -1368
rect -2950 -1448 2949 -1432
rect -2950 -1512 2865 -1448
rect 2929 -1512 2949 -1448
rect -2950 -1528 2949 -1512
rect -2950 -1592 2865 -1528
rect 2929 -1592 2949 -1528
rect -2950 -1608 2949 -1592
rect -2950 -1672 2865 -1608
rect 2929 -1672 2949 -1608
rect -2950 -1688 2949 -1672
rect -2950 -1752 2865 -1688
rect 2929 -1752 2949 -1688
rect -2950 -1768 2949 -1752
rect -2950 -1832 2865 -1768
rect 2929 -1832 2949 -1768
rect -2950 -1848 2949 -1832
rect -2950 -1912 2865 -1848
rect 2929 -1912 2949 -1848
rect -2950 -1928 2949 -1912
rect -2950 -1992 2865 -1928
rect 2929 -1992 2949 -1928
rect -2950 -2008 2949 -1992
rect -2950 -2072 2865 -2008
rect 2929 -2072 2949 -2008
rect -2950 -2088 2949 -2072
rect -2950 -2152 2865 -2088
rect 2929 -2152 2949 -2088
rect -2950 -2168 2949 -2152
rect -2950 -2232 2865 -2168
rect 2929 -2232 2949 -2168
rect -2950 -2248 2949 -2232
rect -2950 -2312 2865 -2248
rect 2929 -2312 2949 -2248
rect -2950 -2328 2949 -2312
rect -2950 -2392 2865 -2328
rect 2929 -2392 2949 -2328
rect -2950 -2408 2949 -2392
rect -2950 -2472 2865 -2408
rect 2929 -2472 2949 -2408
rect -2950 -2488 2949 -2472
rect -2950 -2552 2865 -2488
rect 2929 -2552 2949 -2488
rect -2950 -2568 2949 -2552
rect -2950 -2632 2865 -2568
rect 2929 -2632 2949 -2568
rect -2950 -2648 2949 -2632
rect -2950 -2712 2865 -2648
rect 2929 -2712 2949 -2648
rect -2950 -2728 2949 -2712
rect -2950 -2792 2865 -2728
rect 2929 -2792 2949 -2728
rect -2950 -2808 2949 -2792
rect -2950 -2872 2865 -2808
rect 2929 -2872 2949 -2808
rect -2950 -2900 2949 -2872
<< via3 >>
rect 2865 2808 2929 2872
rect 2865 2728 2929 2792
rect 2865 2648 2929 2712
rect 2865 2568 2929 2632
rect 2865 2488 2929 2552
rect 2865 2408 2929 2472
rect 2865 2328 2929 2392
rect 2865 2248 2929 2312
rect 2865 2168 2929 2232
rect 2865 2088 2929 2152
rect 2865 2008 2929 2072
rect 2865 1928 2929 1992
rect 2865 1848 2929 1912
rect 2865 1768 2929 1832
rect 2865 1688 2929 1752
rect 2865 1608 2929 1672
rect 2865 1528 2929 1592
rect 2865 1448 2929 1512
rect 2865 1368 2929 1432
rect 2865 1288 2929 1352
rect 2865 1208 2929 1272
rect 2865 1128 2929 1192
rect 2865 1048 2929 1112
rect 2865 968 2929 1032
rect 2865 888 2929 952
rect 2865 808 2929 872
rect 2865 728 2929 792
rect 2865 648 2929 712
rect 2865 568 2929 632
rect 2865 488 2929 552
rect 2865 408 2929 472
rect 2865 328 2929 392
rect 2865 248 2929 312
rect 2865 168 2929 232
rect 2865 88 2929 152
rect 2865 8 2929 72
rect 2865 -72 2929 -8
rect 2865 -152 2929 -88
rect 2865 -232 2929 -168
rect 2865 -312 2929 -248
rect 2865 -392 2929 -328
rect 2865 -472 2929 -408
rect 2865 -552 2929 -488
rect 2865 -632 2929 -568
rect 2865 -712 2929 -648
rect 2865 -792 2929 -728
rect 2865 -872 2929 -808
rect 2865 -952 2929 -888
rect 2865 -1032 2929 -968
rect 2865 -1112 2929 -1048
rect 2865 -1192 2929 -1128
rect 2865 -1272 2929 -1208
rect 2865 -1352 2929 -1288
rect 2865 -1432 2929 -1368
rect 2865 -1512 2929 -1448
rect 2865 -1592 2929 -1528
rect 2865 -1672 2929 -1608
rect 2865 -1752 2929 -1688
rect 2865 -1832 2929 -1768
rect 2865 -1912 2929 -1848
rect 2865 -1992 2929 -1928
rect 2865 -2072 2929 -2008
rect 2865 -2152 2929 -2088
rect 2865 -2232 2929 -2168
rect 2865 -2312 2929 -2248
rect 2865 -2392 2929 -2328
rect 2865 -2472 2929 -2408
rect 2865 -2552 2929 -2488
rect 2865 -2632 2929 -2568
rect 2865 -2712 2929 -2648
rect 2865 -2792 2929 -2728
rect 2865 -2872 2929 -2808
<< mimcap >>
rect -2850 2752 2750 2800
rect -2850 -2752 -2802 2752
rect 2702 -2752 2750 2752
rect -2850 -2800 2750 -2752
<< mimcapcontact >>
rect -2802 -2752 2702 2752
<< metal4 >>
rect 2849 2872 2945 2888
rect 2849 2808 2865 2872
rect 2929 2808 2945 2872
rect 2849 2792 2945 2808
rect -2811 2752 2711 2761
rect -2811 -2752 -2802 2752
rect 2702 -2752 2711 2752
rect -2811 -2761 2711 -2752
rect 2849 2728 2865 2792
rect 2929 2728 2945 2792
rect 2849 2712 2945 2728
rect 2849 2648 2865 2712
rect 2929 2648 2945 2712
rect 2849 2632 2945 2648
rect 2849 2568 2865 2632
rect 2929 2568 2945 2632
rect 2849 2552 2945 2568
rect 2849 2488 2865 2552
rect 2929 2488 2945 2552
rect 2849 2472 2945 2488
rect 2849 2408 2865 2472
rect 2929 2408 2945 2472
rect 2849 2392 2945 2408
rect 2849 2328 2865 2392
rect 2929 2328 2945 2392
rect 2849 2312 2945 2328
rect 2849 2248 2865 2312
rect 2929 2248 2945 2312
rect 2849 2232 2945 2248
rect 2849 2168 2865 2232
rect 2929 2168 2945 2232
rect 2849 2152 2945 2168
rect 2849 2088 2865 2152
rect 2929 2088 2945 2152
rect 2849 2072 2945 2088
rect 2849 2008 2865 2072
rect 2929 2008 2945 2072
rect 2849 1992 2945 2008
rect 2849 1928 2865 1992
rect 2929 1928 2945 1992
rect 2849 1912 2945 1928
rect 2849 1848 2865 1912
rect 2929 1848 2945 1912
rect 2849 1832 2945 1848
rect 2849 1768 2865 1832
rect 2929 1768 2945 1832
rect 2849 1752 2945 1768
rect 2849 1688 2865 1752
rect 2929 1688 2945 1752
rect 2849 1672 2945 1688
rect 2849 1608 2865 1672
rect 2929 1608 2945 1672
rect 2849 1592 2945 1608
rect 2849 1528 2865 1592
rect 2929 1528 2945 1592
rect 2849 1512 2945 1528
rect 2849 1448 2865 1512
rect 2929 1448 2945 1512
rect 2849 1432 2945 1448
rect 2849 1368 2865 1432
rect 2929 1368 2945 1432
rect 2849 1352 2945 1368
rect 2849 1288 2865 1352
rect 2929 1288 2945 1352
rect 2849 1272 2945 1288
rect 2849 1208 2865 1272
rect 2929 1208 2945 1272
rect 2849 1192 2945 1208
rect 2849 1128 2865 1192
rect 2929 1128 2945 1192
rect 2849 1112 2945 1128
rect 2849 1048 2865 1112
rect 2929 1048 2945 1112
rect 2849 1032 2945 1048
rect 2849 968 2865 1032
rect 2929 968 2945 1032
rect 2849 952 2945 968
rect 2849 888 2865 952
rect 2929 888 2945 952
rect 2849 872 2945 888
rect 2849 808 2865 872
rect 2929 808 2945 872
rect 2849 792 2945 808
rect 2849 728 2865 792
rect 2929 728 2945 792
rect 2849 712 2945 728
rect 2849 648 2865 712
rect 2929 648 2945 712
rect 2849 632 2945 648
rect 2849 568 2865 632
rect 2929 568 2945 632
rect 2849 552 2945 568
rect 2849 488 2865 552
rect 2929 488 2945 552
rect 2849 472 2945 488
rect 2849 408 2865 472
rect 2929 408 2945 472
rect 2849 392 2945 408
rect 2849 328 2865 392
rect 2929 328 2945 392
rect 2849 312 2945 328
rect 2849 248 2865 312
rect 2929 248 2945 312
rect 2849 232 2945 248
rect 2849 168 2865 232
rect 2929 168 2945 232
rect 2849 152 2945 168
rect 2849 88 2865 152
rect 2929 88 2945 152
rect 2849 72 2945 88
rect 2849 8 2865 72
rect 2929 8 2945 72
rect 2849 -8 2945 8
rect 2849 -72 2865 -8
rect 2929 -72 2945 -8
rect 2849 -88 2945 -72
rect 2849 -152 2865 -88
rect 2929 -152 2945 -88
rect 2849 -168 2945 -152
rect 2849 -232 2865 -168
rect 2929 -232 2945 -168
rect 2849 -248 2945 -232
rect 2849 -312 2865 -248
rect 2929 -312 2945 -248
rect 2849 -328 2945 -312
rect 2849 -392 2865 -328
rect 2929 -392 2945 -328
rect 2849 -408 2945 -392
rect 2849 -472 2865 -408
rect 2929 -472 2945 -408
rect 2849 -488 2945 -472
rect 2849 -552 2865 -488
rect 2929 -552 2945 -488
rect 2849 -568 2945 -552
rect 2849 -632 2865 -568
rect 2929 -632 2945 -568
rect 2849 -648 2945 -632
rect 2849 -712 2865 -648
rect 2929 -712 2945 -648
rect 2849 -728 2945 -712
rect 2849 -792 2865 -728
rect 2929 -792 2945 -728
rect 2849 -808 2945 -792
rect 2849 -872 2865 -808
rect 2929 -872 2945 -808
rect 2849 -888 2945 -872
rect 2849 -952 2865 -888
rect 2929 -952 2945 -888
rect 2849 -968 2945 -952
rect 2849 -1032 2865 -968
rect 2929 -1032 2945 -968
rect 2849 -1048 2945 -1032
rect 2849 -1112 2865 -1048
rect 2929 -1112 2945 -1048
rect 2849 -1128 2945 -1112
rect 2849 -1192 2865 -1128
rect 2929 -1192 2945 -1128
rect 2849 -1208 2945 -1192
rect 2849 -1272 2865 -1208
rect 2929 -1272 2945 -1208
rect 2849 -1288 2945 -1272
rect 2849 -1352 2865 -1288
rect 2929 -1352 2945 -1288
rect 2849 -1368 2945 -1352
rect 2849 -1432 2865 -1368
rect 2929 -1432 2945 -1368
rect 2849 -1448 2945 -1432
rect 2849 -1512 2865 -1448
rect 2929 -1512 2945 -1448
rect 2849 -1528 2945 -1512
rect 2849 -1592 2865 -1528
rect 2929 -1592 2945 -1528
rect 2849 -1608 2945 -1592
rect 2849 -1672 2865 -1608
rect 2929 -1672 2945 -1608
rect 2849 -1688 2945 -1672
rect 2849 -1752 2865 -1688
rect 2929 -1752 2945 -1688
rect 2849 -1768 2945 -1752
rect 2849 -1832 2865 -1768
rect 2929 -1832 2945 -1768
rect 2849 -1848 2945 -1832
rect 2849 -1912 2865 -1848
rect 2929 -1912 2945 -1848
rect 2849 -1928 2945 -1912
rect 2849 -1992 2865 -1928
rect 2929 -1992 2945 -1928
rect 2849 -2008 2945 -1992
rect 2849 -2072 2865 -2008
rect 2929 -2072 2945 -2008
rect 2849 -2088 2945 -2072
rect 2849 -2152 2865 -2088
rect 2929 -2152 2945 -2088
rect 2849 -2168 2945 -2152
rect 2849 -2232 2865 -2168
rect 2929 -2232 2945 -2168
rect 2849 -2248 2945 -2232
rect 2849 -2312 2865 -2248
rect 2929 -2312 2945 -2248
rect 2849 -2328 2945 -2312
rect 2849 -2392 2865 -2328
rect 2929 -2392 2945 -2328
rect 2849 -2408 2945 -2392
rect 2849 -2472 2865 -2408
rect 2929 -2472 2945 -2408
rect 2849 -2488 2945 -2472
rect 2849 -2552 2865 -2488
rect 2929 -2552 2945 -2488
rect 2849 -2568 2945 -2552
rect 2849 -2632 2865 -2568
rect 2929 -2632 2945 -2568
rect 2849 -2648 2945 -2632
rect 2849 -2712 2865 -2648
rect 2929 -2712 2945 -2648
rect 2849 -2728 2945 -2712
rect 2849 -2792 2865 -2728
rect 2929 -2792 2945 -2728
rect 2849 -2808 2945 -2792
rect 2849 -2872 2865 -2808
rect 2929 -2872 2945 -2808
rect 2849 -2888 2945 -2872
<< properties >>
string FIXED_BBOX -2950 -2900 2850 2900
<< end >>
