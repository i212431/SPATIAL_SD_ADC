magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< nwell >>
rect 33364 14450 34170 15442
rect 33364 14365 33685 14450
<< locali >>
rect 34037 15413 34900 15546
rect 34695 14984 34900 15413
rect 34682 14943 34902 14984
rect 34682 14837 34706 14943
rect 34884 14837 34902 14943
rect 34682 14792 34902 14837
<< viali >>
rect 33707 15513 33741 15547
rect 34706 14837 34884 14943
<< metal1 >>
rect 32292 17526 32868 17622
rect 32292 17282 32394 17526
rect 32766 17282 32868 17526
rect 32292 17170 32868 17282
rect 32401 15930 32679 17170
rect 32401 15682 34134 15930
rect 32401 15652 34007 15682
rect 33330 15561 33756 15562
rect 33101 15547 33756 15561
rect 33101 15513 33707 15547
rect 33741 15513 33756 15547
rect 33101 15510 33756 15513
rect 33101 15202 33135 15510
rect 33443 15420 33756 15510
rect 33443 15202 33472 15420
rect 33101 15148 33472 15202
rect 33586 14648 34136 15186
rect 34682 14948 34902 14984
rect 34682 14832 34705 14948
rect 34885 14832 34902 14948
rect 34682 14792 34902 14832
rect 91054 11553 92077 11582
rect 91054 11373 91085 11553
rect 91265 11373 92077 11553
rect 91054 11248 92077 11373
rect 91743 10699 92077 11248
rect 91743 10365 103133 10699
rect 102795 7202 103129 10365
rect 102642 7056 103302 7202
rect 102642 6748 102776 7056
rect 103148 6748 103302 7056
rect 102642 6604 103302 6748
<< via1 >>
rect 32394 17282 32766 17526
rect 33135 15202 33443 15510
rect 34705 14943 34885 14948
rect 34705 14837 34706 14943
rect 34706 14837 34884 14943
rect 34884 14837 34885 14943
rect 34705 14832 34885 14837
rect 91085 11373 91265 11553
rect 102776 6748 103148 7056
<< metal2 >>
rect 33598 18564 36202 18570
rect 32380 17526 32780 17550
rect 32380 17282 32394 17526
rect 32766 17282 32780 17526
rect 32380 17258 32780 17282
rect 33598 17148 33632 18564
rect 36168 17148 36202 18564
rect 33598 17142 36202 17148
rect 49293 16934 60111 18761
rect 99360 16934 114231 18761
rect 149778 16934 166325 18761
rect 130994 16688 139039 16757
rect 85366 16591 85936 16686
rect 85366 16455 85463 16591
rect 85839 16455 85936 16591
rect 85366 16344 85936 16455
rect 33101 15510 33472 15561
rect 33101 15202 33135 15510
rect 33443 15202 33472 15510
rect 33101 15148 33472 15202
rect 35255 15193 35619 15269
rect 34682 14948 34902 14984
rect 34682 14832 34705 14948
rect 34885 14832 34902 14948
rect 34682 14792 34902 14832
rect 35255 14897 35288 15193
rect 35584 14897 35619 15193
rect 35255 14824 35619 14897
rect 85455 14821 85797 16344
rect 130994 16152 131095 16688
rect 131471 16152 139039 16688
rect 130994 16048 139039 16152
rect 138330 14824 139039 16048
rect 153914 15961 154982 16044
rect 153914 15185 154032 15961
rect 154888 15185 154982 15961
rect 184737 15594 189358 16190
rect 184737 15392 185333 15594
rect 153914 15106 154982 15185
rect 183082 15270 185333 15392
rect 39672 14042 40106 14414
rect 27978 12410 30056 12494
rect 27978 11554 28082 12410
rect 29978 11554 30056 12410
rect 27978 11478 30056 11554
rect 91052 11553 91296 11578
rect 91052 11373 91085 11553
rect 91265 11373 91296 11553
rect 91052 11340 91296 11373
rect 154252 9841 154947 15106
rect 183082 14894 183223 15270
rect 183679 14894 185333 15270
rect 183082 14796 185333 14894
rect 188762 14832 189358 15594
rect 29193 9146 59829 9841
rect 59134 5776 59829 9146
rect 73372 5776 74067 9739
rect 81243 9146 112263 9841
rect 102642 7056 103302 7202
rect 102642 7050 102776 7056
rect 103148 7050 103302 7056
rect 102642 6754 102774 7050
rect 103150 6754 103302 7050
rect 102642 6748 102776 6754
rect 103148 6748 103302 6754
rect 102642 6604 103302 6748
rect 59134 5081 74067 5776
rect 111568 6392 112263 9146
rect 111568 5778 120309 6392
rect 124918 5778 125613 9783
rect 132988 9146 163999 9841
rect 111568 5697 125613 5778
rect 119614 5083 125613 5697
rect 163304 5670 163999 9146
rect 176474 5670 177169 9675
rect 163304 4975 177169 5670
rect 48677 2884 63195 4711
rect 98126 2884 115995 4711
rect 153392 2884 167295 4711
<< via2 >>
rect 33632 17148 36168 18564
rect 85463 16455 85839 16591
rect 33141 15208 33437 15504
rect 35288 14897 35584 15193
rect 131095 16152 131471 16688
rect 154032 15185 154888 15961
rect 28082 11554 29978 12410
rect 91107 11395 91243 11531
rect 183223 14894 183679 15270
rect 102774 6754 102776 7050
rect 102776 6754 103148 7050
rect 103148 6754 103150 7050
<< metal3 >>
rect 33378 18564 36400 18768
rect 33378 17148 33632 18564
rect 36168 18523 36400 18564
rect 36178 17179 36400 18523
rect 36168 17148 36400 17179
rect 33378 16944 36400 17148
rect 89462 18054 90868 21832
rect 89462 17270 89943 18054
rect 90487 17270 90868 18054
rect 193208 19859 194056 21630
rect 89462 16808 90868 17270
rect 141568 17343 142606 17430
rect 141568 17039 141658 17343
rect 142522 17039 142606 17343
rect 141568 16948 142606 17039
rect 193208 17235 193301 19859
rect 193925 17235 194056 19859
rect 85366 16595 85920 16686
rect 85366 16451 85459 16595
rect 85843 16451 85920 16595
rect 85366 16344 85920 16451
rect 33101 15508 33472 15561
rect 33101 15204 33137 15508
rect 33441 15204 33472 15508
rect 33101 15148 33472 15204
rect 35255 15197 35619 15269
rect 35255 14893 35285 15197
rect 35589 14893 35619 15197
rect 35255 14824 35619 14893
rect 39672 14412 40106 14414
rect 39670 14342 40106 14412
rect 39670 14154 39735 14342
rect 39672 14118 39735 14154
rect 40039 14118 40106 14342
rect 39672 14042 40106 14118
rect 38304 12534 38870 12604
rect 27978 12410 30056 12494
rect 27978 12374 28082 12410
rect 29978 12374 30056 12410
rect 27978 11590 28078 12374
rect 29982 11590 30056 12374
rect 38304 12310 38355 12534
rect 38819 12310 38870 12534
rect 38304 12236 38870 12310
rect 90098 12232 90550 16808
rect 131018 16692 131541 16751
rect 131018 16148 131091 16692
rect 131475 16148 131541 16692
rect 131018 16098 131541 16148
rect 91494 12821 91784 14436
rect 91007 12531 91784 12821
rect 27978 11554 28082 11590
rect 29978 11554 30056 11590
rect 27978 11478 30056 11554
rect 91007 11531 91297 12531
rect 91494 12400 91784 12531
rect 141932 12409 142159 16948
rect 193208 16942 194056 17235
rect 194704 17072 195292 17180
rect 153914 15965 154982 16044
rect 153914 15181 154028 15965
rect 154892 15181 154982 15965
rect 153914 15106 154982 15181
rect 183106 15270 183820 15368
rect 183106 15234 183223 15270
rect 183679 15234 183820 15270
rect 183106 14930 183219 15234
rect 183683 14930 183820 15234
rect 183106 14894 183223 14930
rect 183679 14894 183820 14930
rect 183106 14796 183820 14894
rect 193606 12340 194006 16942
rect 194704 16484 204850 17072
rect 194704 14236 195292 16484
rect 204262 16340 204850 16484
rect 204262 16135 206072 16340
rect 204262 15191 204472 16135
rect 205896 15191 206072 16135
rect 204262 14986 206072 15191
rect 91007 11395 91107 11531
rect 91243 11395 91297 11531
rect 91007 11341 91297 11395
rect 102642 7054 103302 7202
rect 102642 6750 102770 7054
rect 103154 6750 103302 7054
rect 102642 6604 103302 6750
<< via3 >>
rect 33634 17179 36168 18523
rect 36168 17179 36178 18523
rect 89943 17270 90487 18054
rect 141658 17039 142522 17343
rect 193301 17235 193925 19859
rect 85459 16591 85843 16595
rect 85459 16455 85463 16591
rect 85463 16455 85839 16591
rect 85839 16455 85843 16591
rect 85459 16451 85843 16455
rect 33137 15504 33441 15508
rect 33137 15208 33141 15504
rect 33141 15208 33437 15504
rect 33437 15208 33441 15504
rect 33137 15204 33441 15208
rect 35285 15193 35589 15197
rect 35285 14897 35288 15193
rect 35288 14897 35584 15193
rect 35584 14897 35589 15193
rect 35285 14893 35589 14897
rect 39735 14118 40039 14342
rect 28078 11590 28082 12374
rect 28082 11590 29978 12374
rect 29978 11590 29982 12374
rect 38355 12310 38819 12534
rect 131091 16688 131475 16692
rect 131091 16152 131095 16688
rect 131095 16152 131471 16688
rect 131471 16152 131475 16688
rect 131091 16148 131475 16152
rect 154028 15961 154892 15965
rect 154028 15185 154032 15961
rect 154032 15185 154888 15961
rect 154888 15185 154892 15961
rect 154028 15181 154892 15185
rect 183219 14930 183223 15234
rect 183223 14930 183679 15234
rect 183679 14930 183683 15234
rect 204472 15191 205896 16135
rect 102770 7050 103154 7054
rect 102770 6754 102774 7050
rect 102774 6754 103150 7050
rect 103150 6754 103154 7050
rect 102770 6750 103154 6754
<< metal4 >>
rect 7200 21155 9516 21558
rect 7200 19319 7436 21155
rect 9272 19319 9516 21155
rect 7200 19074 9516 19319
rect 89462 19704 90868 21832
rect 33378 18523 36390 18758
rect 33378 17179 33634 18523
rect 36178 17179 36390 18523
rect 33378 16932 36390 17179
rect 89462 17228 89752 19704
rect 90628 17228 90868 19704
rect 89462 16808 90868 17228
rect 141568 17343 142612 21648
rect 141568 17309 141658 17343
rect 142522 17309 142612 17343
rect 141568 17073 141652 17309
rect 142528 17073 142612 17309
rect 141568 17039 141658 17073
rect 142522 17039 142612 17073
rect 141568 16942 142612 17039
rect 193208 19859 194056 21630
rect 193208 17235 193301 19859
rect 193925 17235 194056 19859
rect 193208 16942 194056 17235
rect 131159 16751 162009 16756
rect 131018 16692 162009 16751
rect 85366 16595 85920 16686
rect 85366 16451 85459 16595
rect 85843 16451 85920 16595
rect 85366 16447 85920 16451
rect 79691 16338 110038 16447
rect 33101 15508 33472 15561
rect 33101 15204 33137 15508
rect 33441 15204 33472 15508
rect 33101 15148 33472 15204
rect 35254 15280 35642 15282
rect 35254 15197 58476 15280
rect 35254 15174 35285 15197
rect 35256 14893 35285 15174
rect 35589 15171 58476 15197
rect 35589 14893 35619 15171
rect 35256 14824 35619 14893
rect 58367 14966 58476 15171
rect 58367 14857 61717 14966
rect 39672 14412 40106 14414
rect 39670 14348 40106 14412
rect 39670 14342 39769 14348
rect 40005 14342 40106 14348
rect 39670 14154 39735 14342
rect 39672 14118 39735 14154
rect 40039 14118 40106 14342
rect 61608 14330 61717 14857
rect 79691 14802 79800 16338
rect 72458 14693 79800 14802
rect 80485 15825 109121 16147
rect 72458 14330 72567 14693
rect 80485 14465 80807 15825
rect 61608 14221 72567 14330
rect 39672 14112 39769 14118
rect 40005 14112 40106 14118
rect 39672 14042 40106 14112
rect 72743 14143 80807 14465
rect 49350 13808 51238 13960
rect 49350 13755 49531 13808
rect 44165 13572 49531 13755
rect 49767 13572 49851 13808
rect 50087 13572 50171 13808
rect 50407 13572 50491 13808
rect 50727 13572 50811 13808
rect 51047 13755 51238 13808
rect 72743 13755 73065 14143
rect 51047 13572 73065 13755
rect 44165 13433 73065 13572
rect 93220 13712 93616 13770
rect 93220 13476 93301 13712
rect 93537 13476 93616 13712
rect 93220 13420 93616 13476
rect 96183 13389 96505 15825
rect 108799 13207 109121 15825
rect 109929 13671 110038 16338
rect 131018 16148 131091 16692
rect 131475 16647 162009 16692
rect 131475 16148 131541 16647
rect 131018 16098 131541 16148
rect 131957 16427 148319 16433
rect 131957 16111 153289 16427
rect 131159 14911 131268 16098
rect 122700 14802 131268 14911
rect 122700 13671 122809 14802
rect 131957 14535 132279 16111
rect 147997 16105 153289 16111
rect 109929 13562 122809 13671
rect 123415 14213 132279 14535
rect 143170 14484 143626 14544
rect 143170 14248 143287 14484
rect 143523 14248 143626 14484
rect 123415 13207 123737 14213
rect 143170 14174 143626 14248
rect 144892 13743 145442 13800
rect 144892 13507 145054 13743
rect 145290 13507 145442 13743
rect 144892 13420 145442 13507
rect 147997 13489 148319 16105
rect 152967 14573 153289 16105
rect 153914 15965 154982 16044
rect 153914 15851 154028 15965
rect 154892 15851 154982 15965
rect 153914 15295 154022 15851
rect 154898 15295 154982 15851
rect 153914 15181 154028 15295
rect 154892 15181 154982 15295
rect 153914 15106 154982 15181
rect 161900 14899 162009 16647
rect 184063 16367 200489 16689
rect 183106 15234 183820 15368
rect 183106 14930 183219 15234
rect 183683 14930 183820 15234
rect 183106 14899 183820 14930
rect 161900 14796 183820 14899
rect 161900 14790 183779 14796
rect 184063 14573 184385 16367
rect 152967 14251 184385 14573
rect 196680 13723 197182 13860
rect 196680 13487 196812 13723
rect 197048 13487 197182 13723
rect 200167 13557 200489 16367
rect 204278 16135 206056 16326
rect 204278 15191 204472 16135
rect 205896 15191 206056 16135
rect 204278 15000 206056 15191
rect 196680 13358 197182 13487
rect 108799 12885 123737 13207
rect 38304 12540 38870 12604
rect 38304 12534 38469 12540
rect 38705 12534 38870 12540
rect 27978 12374 30056 12494
rect 27978 11590 28078 12374
rect 29982 11590 30056 12374
rect 38304 12310 38355 12534
rect 38819 12310 38870 12534
rect 38304 12304 38469 12310
rect 38705 12304 38870 12310
rect 38304 12236 38870 12304
rect 153716 12168 154386 12270
rect 102090 11908 102523 12009
rect 27978 11478 30056 11590
rect 50342 11710 50972 11856
rect 50342 11474 50631 11710
rect 50867 11474 50972 11710
rect 102090 11672 102209 11908
rect 102445 11672 102523 11908
rect 102090 11576 102523 11672
rect 153716 11932 153927 12168
rect 154163 11932 154386 12168
rect 153716 11502 154386 11932
rect 50342 11390 50972 11474
rect 102642 7054 103302 7202
rect 102642 6750 102770 7054
rect 103154 6750 103302 7054
rect 102642 6604 103302 6750
<< via4 >>
rect 7436 19319 9272 21155
rect 33668 17253 36144 18449
rect 89752 18054 90628 19704
rect 89752 17270 89943 18054
rect 89943 17270 90487 18054
rect 90487 17270 90628 18054
rect 89752 17228 90628 17270
rect 141652 17073 141658 17309
rect 141658 17073 141888 17309
rect 141972 17073 142208 17309
rect 142292 17073 142522 17309
rect 142522 17073 142528 17309
rect 193335 17309 193891 19785
rect 33171 15238 33407 15474
rect 39769 14342 40005 14348
rect 39769 14118 40005 14342
rect 39769 14112 40005 14118
rect 49531 13572 49767 13808
rect 49851 13572 50087 13808
rect 50171 13572 50407 13808
rect 50491 13572 50727 13808
rect 50811 13572 51047 13808
rect 93301 13476 93537 13712
rect 143287 14248 143523 14484
rect 145054 13507 145290 13743
rect 154022 15295 154028 15851
rect 154028 15295 154892 15851
rect 154892 15295 154898 15851
rect 196812 13487 197048 13723
rect 204586 15225 205782 16101
rect 38469 12534 38705 12540
rect 28112 11704 29948 12260
rect 38469 12310 38705 12534
rect 38469 12304 38705 12310
rect 50631 11474 50867 11710
rect 102209 11672 102445 11908
rect 153927 11932 154163 12168
rect 102844 6784 103080 7020
<< metal5 >>
rect 7200 21155 9516 21558
rect 7200 19319 7436 21155
rect 9272 19319 9516 21155
rect 7200 19074 9516 19319
rect 33376 18449 36396 21772
rect 33376 17253 33668 18449
rect 36144 17253 36396 18449
rect 33376 16940 36396 17253
rect 42030 16683 43057 21733
rect 38297 16117 43057 16683
rect 38304 15845 43057 16117
rect 32972 15627 33523 15629
rect 20321 15474 33523 15627
rect 20321 15238 33171 15474
rect 33407 15238 33523 15474
rect 20321 15122 33523 15238
rect 20321 3437 20826 15122
rect 32972 15106 33523 15122
rect 38304 12540 38870 15845
rect 27970 12260 30056 12496
rect 27970 11704 28112 12260
rect 29948 11704 30056 12260
rect 38304 12304 38469 12540
rect 38705 12304 38870 12540
rect 38304 12236 38870 12304
rect 39672 14348 40106 14414
rect 39672 14112 39769 14348
rect 40005 14112 40106 14348
rect 39672 11797 40106 14112
rect 49350 13808 51240 21634
rect 89462 19704 90868 21832
rect 89462 17228 89752 19704
rect 90628 17228 90868 19704
rect 89462 16808 90868 17228
rect 141568 17309 142612 21648
rect 141568 17073 141652 17309
rect 141888 17073 141972 17309
rect 142208 17073 142292 17309
rect 142528 17073 142612 17309
rect 141568 16942 142612 17073
rect 153914 15851 154982 21554
rect 193208 19785 194056 21630
rect 193208 17309 193335 19785
rect 193891 17309 194056 19785
rect 193208 16942 194056 17309
rect 153914 15295 154022 15851
rect 154898 15295 154982 15851
rect 153914 15104 154982 15295
rect 204244 16101 206056 16326
rect 204244 15225 204586 16101
rect 205782 15225 206056 16101
rect 143168 14484 146512 14544
rect 143168 14248 143287 14484
rect 143523 14248 146512 14484
rect 143168 14176 146512 14248
rect 143170 14174 143626 14176
rect 93006 13811 93612 13902
rect 146062 13888 146512 14176
rect 49350 13572 49531 13808
rect 49767 13572 49851 13808
rect 50087 13572 50171 13808
rect 50407 13572 50491 13808
rect 50727 13572 50811 13808
rect 51047 13572 51240 13808
rect 49350 13434 51240 13572
rect 53216 13712 93636 13811
rect 53216 13476 93301 13712
rect 93537 13476 93636 13712
rect 53216 13378 93636 13476
rect 144904 13743 145554 13798
rect 144904 13507 145054 13743
rect 145290 13507 145554 13743
rect 27970 11480 30056 11704
rect 36905 11363 40106 11797
rect 50342 11823 50972 11856
rect 53216 11823 53649 13378
rect 144904 12756 145554 13507
rect 146062 13438 151501 13888
rect 144876 12371 145554 12756
rect 50342 11710 53649 11823
rect 50342 11474 50631 11710
rect 50867 11474 53649 11710
rect 102090 12323 145554 12371
rect 102090 11938 145534 12323
rect 102090 11908 102523 11938
rect 102090 11672 102209 11908
rect 102445 11672 102523 11908
rect 102090 11576 102523 11672
rect 50342 11390 53649 11474
rect 11579 2615 20826 3437
rect 22786 10953 27583 11200
rect 36906 10953 37339 11363
rect 22786 10520 37339 10953
rect 11579 -199 12508 2615
rect 22786 -112 23545 10520
rect 102482 7020 103640 7222
rect 102482 6784 102844 7020
rect 103080 6784 103640 7020
rect 102482 -304 103640 6784
rect 151051 -157 151501 13438
rect 196677 13723 198308 14113
rect 196677 13487 196812 13723
rect 197048 13487 198308 13723
rect 196677 13343 198308 13487
rect 197538 12268 198308 13343
rect 153720 12168 198308 12268
rect 153720 11932 153927 12168
rect 154163 11932 198308 12168
rect 153720 11498 198308 11932
rect 204244 -546 206056 15225
use TOP1nn  TOP1nn_0
timestamp 1667803582
transform 1 0 30608 0 1 13484
box -30608 -13484 25640 8020
use TOP2nn  TOP2nn_0
timestamp 1667803582
transform 1 0 82366 0 1 13484
box -30608 -13484 25640 8020
use TOP2nn  TOP2nn_1
timestamp 1667803582
transform 1 0 134111 0 1 13484
box -30608 -13484 25640 8020
use TOP2nn  TOP2nn_2
timestamp 1667803582
transform 1 0 185873 0 1 13484
box -30608 -13484 25640 8020
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_0
timestamp 1667803582
transform 1 0 33586 0 -1 15700
box -38 -48 590 592
<< labels >>
flabel metal5 s 154452 21516 154452 21516 0 FreeSans 16000 0 0 0 IBIAS
port 1 nsew
flabel metal5 s 8282 21520 8282 21520 0 FreeSans 16000 0 0 0 VSS
port 2 nsew
flabel metal5 s 34782 21524 34782 21524 0 FreeSans 16000 0 0 0 VDD
port 3 nsew
flabel metal5 s 50180 21594 50180 21594 0 FreeSans 16000 0 0 0 VREF
port 4 nsew
flabel metal5 s 42774 21616 42774 21616 0 FreeSans 14000 0 0 0 SD_IN_1
port 5 nsew
flabel metal5 s 23328 -82 23328 -82 0 FreeSans 16000 0 0 0 SD_DOUT_1
port 6 nsew
flabel metal5 s 102924 -74 102924 -74 0 FreeSans 16000 0 0 0 SD_DOUT_2
port 7 nsew
flabel metal5 s 89904 21634 89904 21634 0 FreeSans 16000 0 0 0 SD_IN_2
port 8 nsew
flabel metal5 s 142044 21590 142044 21590 0 FreeSans 16000 0 0 0 SD_IN_3
port 9 nsew
flabel metal5 s 151276 -58 151276 -58 0 FreeSans 16000 0 0 0 SD_DOUT_3
port 10 nsew
flabel metal5 s 193626 21584 193626 21584 0 FreeSans 16000 0 0 0 SD_IN_4
port 11 nsew
flabel metal5 s 205038 -268 205038 -268 0 FreeSans 16000 0 0 0 SD_DOUT_4
port 12 nsew
flabel metal5 s 12249 -89 12249 -89 0 FreeSans 16000 0 0 0 CLK
port 13 nsew
<< end >>
