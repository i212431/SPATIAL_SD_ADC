magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< error_p >>
rect -77 322 -19 328
rect 115 322 173 328
rect -77 288 -65 322
rect 115 288 127 322
rect -77 282 -19 288
rect 115 282 173 288
rect -173 -288 -115 -282
rect 19 -288 77 -282
rect -173 -322 -161 -288
rect 19 -322 31 -288
rect -173 -328 -115 -322
rect 19 -328 77 -322
<< pwell >>
rect -247 -276 247 276
<< nmos >>
rect -159 -250 -129 250
rect -63 -250 -33 250
rect 33 -250 63 250
rect 129 -250 159 250
<< ndiff >>
rect -221 221 -159 250
rect -221 187 -209 221
rect -175 187 -159 221
rect -221 153 -159 187
rect -221 119 -209 153
rect -175 119 -159 153
rect -221 85 -159 119
rect -221 51 -209 85
rect -175 51 -159 85
rect -221 17 -159 51
rect -221 -17 -209 17
rect -175 -17 -159 17
rect -221 -51 -159 -17
rect -221 -85 -209 -51
rect -175 -85 -159 -51
rect -221 -119 -159 -85
rect -221 -153 -209 -119
rect -175 -153 -159 -119
rect -221 -187 -159 -153
rect -221 -221 -209 -187
rect -175 -221 -159 -187
rect -221 -250 -159 -221
rect -129 221 -63 250
rect -129 187 -113 221
rect -79 187 -63 221
rect -129 153 -63 187
rect -129 119 -113 153
rect -79 119 -63 153
rect -129 85 -63 119
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -119 -63 -85
rect -129 -153 -113 -119
rect -79 -153 -63 -119
rect -129 -187 -63 -153
rect -129 -221 -113 -187
rect -79 -221 -63 -187
rect -129 -250 -63 -221
rect -33 221 33 250
rect -33 187 -17 221
rect 17 187 33 221
rect -33 153 33 187
rect -33 119 -17 153
rect 17 119 33 153
rect -33 85 33 119
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -119 33 -85
rect -33 -153 -17 -119
rect 17 -153 33 -119
rect -33 -187 33 -153
rect -33 -221 -17 -187
rect 17 -221 33 -187
rect -33 -250 33 -221
rect 63 221 129 250
rect 63 187 79 221
rect 113 187 129 221
rect 63 153 129 187
rect 63 119 79 153
rect 113 119 129 153
rect 63 85 129 119
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -119 129 -85
rect 63 -153 79 -119
rect 113 -153 129 -119
rect 63 -187 129 -153
rect 63 -221 79 -187
rect 113 -221 129 -187
rect 63 -250 129 -221
rect 159 221 221 250
rect 159 187 175 221
rect 209 187 221 221
rect 159 153 221 187
rect 159 119 175 153
rect 209 119 221 153
rect 159 85 221 119
rect 159 51 175 85
rect 209 51 221 85
rect 159 17 221 51
rect 159 -17 175 17
rect 209 -17 221 17
rect 159 -51 221 -17
rect 159 -85 175 -51
rect 209 -85 221 -51
rect 159 -119 221 -85
rect 159 -153 175 -119
rect 209 -153 221 -119
rect 159 -187 221 -153
rect 159 -221 175 -187
rect 209 -221 221 -187
rect 159 -250 221 -221
<< ndiffc >>
rect -209 187 -175 221
rect -209 119 -175 153
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -209 -153 -175 -119
rect -209 -221 -175 -187
rect -113 187 -79 221
rect -113 119 -79 153
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -113 -153 -79 -119
rect -113 -221 -79 -187
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect 79 187 113 221
rect 79 119 113 153
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 79 -153 113 -119
rect 79 -221 113 -187
rect 175 187 209 221
rect 175 119 209 153
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 175 -153 209 -119
rect 175 -221 209 -187
<< poly >>
rect -81 322 -15 338
rect -81 288 -65 322
rect -31 288 -15 322
rect -159 250 -129 276
rect -81 272 -15 288
rect 111 322 177 338
rect 111 288 127 322
rect 161 288 177 322
rect -63 250 -33 272
rect 33 250 63 276
rect 111 272 177 288
rect 129 250 159 272
rect -159 -272 -129 -250
rect -177 -288 -111 -272
rect -63 -276 -33 -250
rect 33 -272 63 -250
rect -177 -322 -161 -288
rect -127 -322 -111 -288
rect -177 -338 -111 -322
rect 15 -288 81 -272
rect 129 -276 159 -250
rect 15 -322 31 -288
rect 65 -322 81 -288
rect 15 -338 81 -322
<< polycont >>
rect -65 288 -31 322
rect 127 288 161 322
rect -161 -322 -127 -288
rect 31 -322 65 -288
<< locali >>
rect -81 288 -65 322
rect -31 288 -15 322
rect 111 288 127 322
rect 161 288 177 322
rect -209 233 -175 254
rect -209 161 -175 187
rect -209 89 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -89
rect -209 -187 -175 -161
rect -209 -254 -175 -233
rect -113 233 -79 254
rect -113 161 -79 187
rect -113 89 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -89
rect -113 -187 -79 -161
rect -113 -254 -79 -233
rect -17 233 17 254
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -254 17 -233
rect 79 233 113 254
rect 79 161 113 187
rect 79 89 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -89
rect 79 -187 113 -161
rect 79 -254 113 -233
rect 175 233 209 254
rect 175 161 209 187
rect 175 89 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -89
rect 175 -187 209 -161
rect 175 -254 209 -233
rect -177 -322 -161 -288
rect -127 -322 -111 -288
rect 15 -322 31 -288
rect 65 -322 81 -288
<< viali >>
rect -65 288 -31 322
rect 127 288 161 322
rect -209 221 -175 233
rect -209 199 -175 221
rect -209 153 -175 161
rect -209 127 -175 153
rect -209 85 -175 89
rect -209 55 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -55
rect -209 -89 -175 -85
rect -209 -153 -175 -127
rect -209 -161 -175 -153
rect -209 -221 -175 -199
rect -209 -233 -175 -221
rect -113 221 -79 233
rect -113 199 -79 221
rect -113 153 -79 161
rect -113 127 -79 153
rect -113 85 -79 89
rect -113 55 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -55
rect -113 -89 -79 -85
rect -113 -153 -79 -127
rect -113 -161 -79 -153
rect -113 -221 -79 -199
rect -113 -233 -79 -221
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect 79 221 113 233
rect 79 199 113 221
rect 79 153 113 161
rect 79 127 113 153
rect 79 85 113 89
rect 79 55 113 85
rect 79 -17 113 17
rect 79 -85 113 -55
rect 79 -89 113 -85
rect 79 -153 113 -127
rect 79 -161 113 -153
rect 79 -221 113 -199
rect 79 -233 113 -221
rect 175 221 209 233
rect 175 199 209 221
rect 175 153 209 161
rect 175 127 209 153
rect 175 85 209 89
rect 175 55 209 85
rect 175 -17 209 17
rect 175 -85 209 -55
rect 175 -89 209 -85
rect 175 -153 209 -127
rect 175 -161 209 -153
rect 175 -221 209 -199
rect 175 -233 209 -221
rect -161 -322 -127 -288
rect 31 -322 65 -288
<< metal1 >>
rect -77 322 -19 328
rect -77 288 -65 322
rect -31 288 -19 322
rect -77 282 -19 288
rect 115 322 173 328
rect 115 288 127 322
rect 161 288 173 322
rect 115 282 173 288
rect -215 233 -169 250
rect -215 199 -209 233
rect -175 199 -169 233
rect -215 161 -169 199
rect -215 127 -209 161
rect -175 127 -169 161
rect -215 89 -169 127
rect -215 55 -209 89
rect -175 55 -169 89
rect -215 17 -169 55
rect -215 -17 -209 17
rect -175 -17 -169 17
rect -215 -55 -169 -17
rect -215 -89 -209 -55
rect -175 -89 -169 -55
rect -215 -127 -169 -89
rect -215 -161 -209 -127
rect -175 -161 -169 -127
rect -215 -199 -169 -161
rect -215 -233 -209 -199
rect -175 -233 -169 -199
rect -215 -250 -169 -233
rect -119 233 -73 250
rect -119 199 -113 233
rect -79 199 -73 233
rect -119 161 -73 199
rect -119 127 -113 161
rect -79 127 -73 161
rect -119 89 -73 127
rect -119 55 -113 89
rect -79 55 -73 89
rect -119 17 -73 55
rect -119 -17 -113 17
rect -79 -17 -73 17
rect -119 -55 -73 -17
rect -119 -89 -113 -55
rect -79 -89 -73 -55
rect -119 -127 -73 -89
rect -119 -161 -113 -127
rect -79 -161 -73 -127
rect -119 -199 -73 -161
rect -119 -233 -113 -199
rect -79 -233 -73 -199
rect -119 -250 -73 -233
rect -23 233 23 250
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -250 23 -233
rect 73 233 119 250
rect 73 199 79 233
rect 113 199 119 233
rect 73 161 119 199
rect 73 127 79 161
rect 113 127 119 161
rect 73 89 119 127
rect 73 55 79 89
rect 113 55 119 89
rect 73 17 119 55
rect 73 -17 79 17
rect 113 -17 119 17
rect 73 -55 119 -17
rect 73 -89 79 -55
rect 113 -89 119 -55
rect 73 -127 119 -89
rect 73 -161 79 -127
rect 113 -161 119 -127
rect 73 -199 119 -161
rect 73 -233 79 -199
rect 113 -233 119 -199
rect 73 -250 119 -233
rect 169 233 215 250
rect 169 199 175 233
rect 209 199 215 233
rect 169 161 215 199
rect 169 127 175 161
rect 209 127 215 161
rect 169 89 215 127
rect 169 55 175 89
rect 209 55 215 89
rect 169 17 215 55
rect 169 -17 175 17
rect 209 -17 215 17
rect 169 -55 215 -17
rect 169 -89 175 -55
rect 209 -89 215 -55
rect 169 -127 215 -89
rect 169 -161 175 -127
rect 209 -161 215 -127
rect 169 -199 215 -161
rect 169 -233 175 -199
rect 209 -233 215 -199
rect 169 -250 215 -233
rect -173 -288 -115 -282
rect -173 -322 -161 -288
rect -127 -322 -115 -288
rect -173 -328 -115 -322
rect 19 -288 77 -282
rect 19 -322 31 -288
rect 65 -322 77 -288
rect 19 -328 77 -322
<< end >>
