magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< error_p >>
rect -77 581 -19 587
rect 115 581 173 587
rect -77 547 -65 581
rect 115 547 127 581
rect -77 541 -19 547
rect 115 541 173 547
rect -173 -547 -115 -541
rect 19 -547 77 -541
rect -173 -581 -161 -547
rect 19 -581 31 -547
rect -173 -587 -115 -581
rect 19 -587 77 -581
<< nwell >>
rect -161 562 257 600
rect -257 -562 257 562
rect -257 -600 161 -562
<< pmos >>
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
<< pdiff >>
rect -221 459 -159 500
rect -221 425 -209 459
rect -175 425 -159 459
rect -221 391 -159 425
rect -221 357 -209 391
rect -175 357 -159 391
rect -221 323 -159 357
rect -221 289 -209 323
rect -175 289 -159 323
rect -221 255 -159 289
rect -221 221 -209 255
rect -175 221 -159 255
rect -221 187 -159 221
rect -221 153 -209 187
rect -175 153 -159 187
rect -221 119 -159 153
rect -221 85 -209 119
rect -175 85 -159 119
rect -221 51 -159 85
rect -221 17 -209 51
rect -175 17 -159 51
rect -221 -17 -159 17
rect -221 -51 -209 -17
rect -175 -51 -159 -17
rect -221 -85 -159 -51
rect -221 -119 -209 -85
rect -175 -119 -159 -85
rect -221 -153 -159 -119
rect -221 -187 -209 -153
rect -175 -187 -159 -153
rect -221 -221 -159 -187
rect -221 -255 -209 -221
rect -175 -255 -159 -221
rect -221 -289 -159 -255
rect -221 -323 -209 -289
rect -175 -323 -159 -289
rect -221 -357 -159 -323
rect -221 -391 -209 -357
rect -175 -391 -159 -357
rect -221 -425 -159 -391
rect -221 -459 -209 -425
rect -175 -459 -159 -425
rect -221 -500 -159 -459
rect -129 459 -63 500
rect -129 425 -113 459
rect -79 425 -63 459
rect -129 391 -63 425
rect -129 357 -113 391
rect -79 357 -63 391
rect -129 323 -63 357
rect -129 289 -113 323
rect -79 289 -63 323
rect -129 255 -63 289
rect -129 221 -113 255
rect -79 221 -63 255
rect -129 187 -63 221
rect -129 153 -113 187
rect -79 153 -63 187
rect -129 119 -63 153
rect -129 85 -113 119
rect -79 85 -63 119
rect -129 51 -63 85
rect -129 17 -113 51
rect -79 17 -63 51
rect -129 -17 -63 17
rect -129 -51 -113 -17
rect -79 -51 -63 -17
rect -129 -85 -63 -51
rect -129 -119 -113 -85
rect -79 -119 -63 -85
rect -129 -153 -63 -119
rect -129 -187 -113 -153
rect -79 -187 -63 -153
rect -129 -221 -63 -187
rect -129 -255 -113 -221
rect -79 -255 -63 -221
rect -129 -289 -63 -255
rect -129 -323 -113 -289
rect -79 -323 -63 -289
rect -129 -357 -63 -323
rect -129 -391 -113 -357
rect -79 -391 -63 -357
rect -129 -425 -63 -391
rect -129 -459 -113 -425
rect -79 -459 -63 -425
rect -129 -500 -63 -459
rect -33 459 33 500
rect -33 425 -17 459
rect 17 425 33 459
rect -33 391 33 425
rect -33 357 -17 391
rect 17 357 33 391
rect -33 323 33 357
rect -33 289 -17 323
rect 17 289 33 323
rect -33 255 33 289
rect -33 221 -17 255
rect 17 221 33 255
rect -33 187 33 221
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -221 33 -187
rect -33 -255 -17 -221
rect 17 -255 33 -221
rect -33 -289 33 -255
rect -33 -323 -17 -289
rect 17 -323 33 -289
rect -33 -357 33 -323
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -33 -425 33 -391
rect -33 -459 -17 -425
rect 17 -459 33 -425
rect -33 -500 33 -459
rect 63 459 129 500
rect 63 425 79 459
rect 113 425 129 459
rect 63 391 129 425
rect 63 357 79 391
rect 113 357 129 391
rect 63 323 129 357
rect 63 289 79 323
rect 113 289 129 323
rect 63 255 129 289
rect 63 221 79 255
rect 113 221 129 255
rect 63 187 129 221
rect 63 153 79 187
rect 113 153 129 187
rect 63 119 129 153
rect 63 85 79 119
rect 113 85 129 119
rect 63 51 129 85
rect 63 17 79 51
rect 113 17 129 51
rect 63 -17 129 17
rect 63 -51 79 -17
rect 113 -51 129 -17
rect 63 -85 129 -51
rect 63 -119 79 -85
rect 113 -119 129 -85
rect 63 -153 129 -119
rect 63 -187 79 -153
rect 113 -187 129 -153
rect 63 -221 129 -187
rect 63 -255 79 -221
rect 113 -255 129 -221
rect 63 -289 129 -255
rect 63 -323 79 -289
rect 113 -323 129 -289
rect 63 -357 129 -323
rect 63 -391 79 -357
rect 113 -391 129 -357
rect 63 -425 129 -391
rect 63 -459 79 -425
rect 113 -459 129 -425
rect 63 -500 129 -459
rect 159 459 221 500
rect 159 425 175 459
rect 209 425 221 459
rect 159 391 221 425
rect 159 357 175 391
rect 209 357 221 391
rect 159 323 221 357
rect 159 289 175 323
rect 209 289 221 323
rect 159 255 221 289
rect 159 221 175 255
rect 209 221 221 255
rect 159 187 221 221
rect 159 153 175 187
rect 209 153 221 187
rect 159 119 221 153
rect 159 85 175 119
rect 209 85 221 119
rect 159 51 221 85
rect 159 17 175 51
rect 209 17 221 51
rect 159 -17 221 17
rect 159 -51 175 -17
rect 209 -51 221 -17
rect 159 -85 221 -51
rect 159 -119 175 -85
rect 209 -119 221 -85
rect 159 -153 221 -119
rect 159 -187 175 -153
rect 209 -187 221 -153
rect 159 -221 221 -187
rect 159 -255 175 -221
rect 209 -255 221 -221
rect 159 -289 221 -255
rect 159 -323 175 -289
rect 209 -323 221 -289
rect 159 -357 221 -323
rect 159 -391 175 -357
rect 209 -391 221 -357
rect 159 -425 221 -391
rect 159 -459 175 -425
rect 209 -459 221 -425
rect 159 -500 221 -459
<< pdiffc >>
rect -209 425 -175 459
rect -209 357 -175 391
rect -209 289 -175 323
rect -209 221 -175 255
rect -209 153 -175 187
rect -209 85 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -85
rect -209 -187 -175 -153
rect -209 -255 -175 -221
rect -209 -323 -175 -289
rect -209 -391 -175 -357
rect -209 -459 -175 -425
rect -113 425 -79 459
rect -113 357 -79 391
rect -113 289 -79 323
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -113 -323 -79 -289
rect -113 -391 -79 -357
rect -113 -459 -79 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 79 425 113 459
rect 79 357 113 391
rect 79 289 113 323
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 79 -323 113 -289
rect 79 -391 113 -357
rect 79 -459 113 -425
rect 175 425 209 459
rect 175 357 209 391
rect 175 289 209 323
rect 175 221 209 255
rect 175 153 209 187
rect 175 85 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -85
rect 175 -187 209 -153
rect 175 -255 209 -221
rect 175 -323 209 -289
rect 175 -391 209 -357
rect 175 -459 209 -425
<< poly >>
rect -81 581 -15 597
rect -81 547 -65 581
rect -31 547 -15 581
rect -81 531 -15 547
rect 111 581 177 597
rect 111 547 127 581
rect 161 547 177 581
rect 111 531 177 547
rect -159 500 -129 526
rect -63 500 -33 531
rect 33 500 63 526
rect 129 500 159 531
rect -159 -531 -129 -500
rect -63 -526 -33 -500
rect 33 -531 63 -500
rect 129 -526 159 -500
rect -177 -547 -111 -531
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect -177 -597 -111 -581
rect 15 -547 81 -531
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 15 -597 81 -581
<< polycont >>
rect -65 547 -31 581
rect 127 547 161 581
rect -161 -581 -127 -547
rect 31 -581 65 -547
<< locali >>
rect -81 547 -65 581
rect -31 547 -15 581
rect 111 547 127 581
rect 161 547 177 581
rect -209 485 -175 504
rect -209 413 -175 425
rect -209 341 -175 357
rect -209 269 -175 289
rect -209 197 -175 221
rect -209 125 -175 153
rect -209 53 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -53
rect -209 -153 -175 -125
rect -209 -221 -175 -197
rect -209 -289 -175 -269
rect -209 -357 -175 -341
rect -209 -425 -175 -413
rect -209 -504 -175 -485
rect -113 485 -79 504
rect -113 413 -79 425
rect -113 341 -79 357
rect -113 269 -79 289
rect -113 197 -79 221
rect -113 125 -79 153
rect -113 53 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -53
rect -113 -153 -79 -125
rect -113 -221 -79 -197
rect -113 -289 -79 -269
rect -113 -357 -79 -341
rect -113 -425 -79 -413
rect -113 -504 -79 -485
rect -17 485 17 504
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -504 17 -485
rect 79 485 113 504
rect 79 413 113 425
rect 79 341 113 357
rect 79 269 113 289
rect 79 197 113 221
rect 79 125 113 153
rect 79 53 113 85
rect 79 -17 113 17
rect 79 -85 113 -53
rect 79 -153 113 -125
rect 79 -221 113 -197
rect 79 -289 113 -269
rect 79 -357 113 -341
rect 79 -425 113 -413
rect 79 -504 113 -485
rect 175 485 209 504
rect 175 413 209 425
rect 175 341 209 357
rect 175 269 209 289
rect 175 197 209 221
rect 175 125 209 153
rect 175 53 209 85
rect 175 -17 209 17
rect 175 -85 209 -53
rect 175 -153 209 -125
rect 175 -221 209 -197
rect 175 -289 209 -269
rect 175 -357 209 -341
rect 175 -425 209 -413
rect 175 -504 209 -485
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect 15 -581 31 -547
rect 65 -581 81 -547
<< viali >>
rect -65 547 -31 581
rect 127 547 161 581
rect -209 459 -175 485
rect -209 451 -175 459
rect -209 391 -175 413
rect -209 379 -175 391
rect -209 323 -175 341
rect -209 307 -175 323
rect -209 255 -175 269
rect -209 235 -175 255
rect -209 187 -175 197
rect -209 163 -175 187
rect -209 119 -175 125
rect -209 91 -175 119
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -209 -119 -175 -91
rect -209 -125 -175 -119
rect -209 -187 -175 -163
rect -209 -197 -175 -187
rect -209 -255 -175 -235
rect -209 -269 -175 -255
rect -209 -323 -175 -307
rect -209 -341 -175 -323
rect -209 -391 -175 -379
rect -209 -413 -175 -391
rect -209 -459 -175 -451
rect -209 -485 -175 -459
rect -113 459 -79 485
rect -113 451 -79 459
rect -113 391 -79 413
rect -113 379 -79 391
rect -113 323 -79 341
rect -113 307 -79 323
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -113 -323 -79 -307
rect -113 -341 -79 -323
rect -113 -391 -79 -379
rect -113 -413 -79 -391
rect -113 -459 -79 -451
rect -113 -485 -79 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 79 459 113 485
rect 79 451 113 459
rect 79 391 113 413
rect 79 379 113 391
rect 79 323 113 341
rect 79 307 113 323
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 79 -323 113 -307
rect 79 -341 113 -323
rect 79 -391 113 -379
rect 79 -413 113 -391
rect 79 -459 113 -451
rect 79 -485 113 -459
rect 175 459 209 485
rect 175 451 209 459
rect 175 391 209 413
rect 175 379 209 391
rect 175 323 209 341
rect 175 307 209 323
rect 175 255 209 269
rect 175 235 209 255
rect 175 187 209 197
rect 175 163 209 187
rect 175 119 209 125
rect 175 91 209 119
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 175 -119 209 -91
rect 175 -125 209 -119
rect 175 -187 209 -163
rect 175 -197 209 -187
rect 175 -255 209 -235
rect 175 -269 209 -255
rect 175 -323 209 -307
rect 175 -341 209 -323
rect 175 -391 209 -379
rect 175 -413 209 -391
rect 175 -459 209 -451
rect 175 -485 209 -459
rect -161 -581 -127 -547
rect 31 -581 65 -547
<< metal1 >>
rect -77 581 -19 587
rect -77 547 -65 581
rect -31 547 -19 581
rect -77 541 -19 547
rect 115 581 173 587
rect 115 547 127 581
rect 161 547 173 581
rect 115 541 173 547
rect -215 485 -169 500
rect -215 451 -209 485
rect -175 451 -169 485
rect -215 413 -169 451
rect -215 379 -209 413
rect -175 379 -169 413
rect -215 341 -169 379
rect -215 307 -209 341
rect -175 307 -169 341
rect -215 269 -169 307
rect -215 235 -209 269
rect -175 235 -169 269
rect -215 197 -169 235
rect -215 163 -209 197
rect -175 163 -169 197
rect -215 125 -169 163
rect -215 91 -209 125
rect -175 91 -169 125
rect -215 53 -169 91
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -91 -169 -53
rect -215 -125 -209 -91
rect -175 -125 -169 -91
rect -215 -163 -169 -125
rect -215 -197 -209 -163
rect -175 -197 -169 -163
rect -215 -235 -169 -197
rect -215 -269 -209 -235
rect -175 -269 -169 -235
rect -215 -307 -169 -269
rect -215 -341 -209 -307
rect -175 -341 -169 -307
rect -215 -379 -169 -341
rect -215 -413 -209 -379
rect -175 -413 -169 -379
rect -215 -451 -169 -413
rect -215 -485 -209 -451
rect -175 -485 -169 -451
rect -215 -500 -169 -485
rect -119 485 -73 500
rect -119 451 -113 485
rect -79 451 -73 485
rect -119 413 -73 451
rect -119 379 -113 413
rect -79 379 -73 413
rect -119 341 -73 379
rect -119 307 -113 341
rect -79 307 -73 341
rect -119 269 -73 307
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -307 -73 -269
rect -119 -341 -113 -307
rect -79 -341 -73 -307
rect -119 -379 -73 -341
rect -119 -413 -113 -379
rect -79 -413 -73 -379
rect -119 -451 -73 -413
rect -119 -485 -113 -451
rect -79 -485 -73 -451
rect -119 -500 -73 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 73 485 119 500
rect 73 451 79 485
rect 113 451 119 485
rect 73 413 119 451
rect 73 379 79 413
rect 113 379 119 413
rect 73 341 119 379
rect 73 307 79 341
rect 113 307 119 341
rect 73 269 119 307
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -307 119 -269
rect 73 -341 79 -307
rect 113 -341 119 -307
rect 73 -379 119 -341
rect 73 -413 79 -379
rect 113 -413 119 -379
rect 73 -451 119 -413
rect 73 -485 79 -451
rect 113 -485 119 -451
rect 73 -500 119 -485
rect 169 485 215 500
rect 169 451 175 485
rect 209 451 215 485
rect 169 413 215 451
rect 169 379 175 413
rect 209 379 215 413
rect 169 341 215 379
rect 169 307 175 341
rect 209 307 215 341
rect 169 269 215 307
rect 169 235 175 269
rect 209 235 215 269
rect 169 197 215 235
rect 169 163 175 197
rect 209 163 215 197
rect 169 125 215 163
rect 169 91 175 125
rect 209 91 215 125
rect 169 53 215 91
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -91 215 -53
rect 169 -125 175 -91
rect 209 -125 215 -91
rect 169 -163 215 -125
rect 169 -197 175 -163
rect 209 -197 215 -163
rect 169 -235 215 -197
rect 169 -269 175 -235
rect 209 -269 215 -235
rect 169 -307 215 -269
rect 169 -341 175 -307
rect 209 -341 215 -307
rect 169 -379 215 -341
rect 169 -413 175 -379
rect 209 -413 215 -379
rect 169 -451 215 -413
rect 169 -485 175 -451
rect 209 -485 215 -451
rect 169 -500 215 -485
rect -173 -547 -115 -541
rect -173 -581 -161 -547
rect -127 -581 -115 -547
rect -173 -587 -115 -581
rect 19 -547 77 -541
rect 19 -581 31 -547
rect 65 -581 77 -547
rect 19 -587 77 -581
<< end >>
