magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< poly >>
rect 41 2408 377 2474
rect 23 1798 360 1864
<< metal1 >>
rect 119 2418 511 2464
rect 70 2336 137 2357
rect 70 2284 77 2336
rect 129 2284 137 2336
rect 70 2262 137 2284
rect 263 2336 329 2357
rect 263 2284 269 2336
rect 321 2284 329 2336
rect 263 2262 329 2284
rect -22 1992 41 2024
rect -22 1940 -17 1992
rect 35 1940 41 1992
rect -22 1907 41 1940
rect 167 1992 233 2024
rect 167 1940 174 1992
rect 226 1940 233 1992
rect 167 1907 233 1940
rect 358 1991 421 2024
rect 358 1939 365 1991
rect 417 1939 421 1991
rect 358 1907 421 1939
rect 465 1854 511 2418
rect 23 1808 511 1854
rect 64 1571 221 1584
rect 64 1519 84 1571
rect 136 1519 148 1571
rect 200 1519 221 1571
rect 64 1507 221 1519
rect 1800 1343 1953 1345
rect 1800 1291 1818 1343
rect 1870 1291 1882 1343
rect 1934 1291 1953 1343
rect 1800 1285 1953 1291
rect 1884 712 2048 719
rect 1884 660 1906 712
rect 1958 660 1970 712
rect 2022 660 2048 712
rect 1884 653 2048 660
rect 65 485 216 497
rect 65 433 82 485
rect 134 433 146 485
rect 198 433 216 485
rect 65 421 216 433
<< via1 >>
rect 77 2284 129 2336
rect 269 2284 321 2336
rect -17 1940 35 1992
rect 174 1940 226 1992
rect 365 1939 417 1991
rect 84 1519 136 1571
rect 148 1519 200 1571
rect 1818 1291 1870 1343
rect 1882 1291 1934 1343
rect 1906 660 1958 712
rect 1970 660 2022 712
rect 82 433 134 485
rect 146 433 198 485
<< metal2 >>
rect 70 2336 600 2357
rect 70 2284 77 2336
rect 129 2284 269 2336
rect 321 2284 600 2336
rect 70 2262 600 2284
rect -32 2023 422 2024
rect -292 1992 422 2023
rect -292 1940 -17 1992
rect 35 1940 174 1992
rect 226 1991 422 1992
rect 226 1940 365 1991
rect -292 1939 365 1940
rect 417 1939 422 1991
rect -292 1916 422 1939
rect -292 1870 -185 1916
rect -32 1907 422 1916
rect -387 1763 -185 1870
rect 54 1571 231 1594
rect 54 1519 84 1571
rect 136 1519 148 1571
rect 200 1519 231 1571
rect 54 485 231 1519
rect 1800 1343 1953 1345
rect 1800 1291 1818 1343
rect 1870 1291 1882 1343
rect 1934 1333 1953 1343
rect 1934 1291 2044 1333
rect 1800 1285 2044 1291
rect 1895 719 2044 1285
rect 2836 735 2984 773
rect 1884 712 2064 719
rect 1884 660 1906 712
rect 1958 660 1970 712
rect 2022 660 2064 712
rect 1884 653 2064 660
rect 2836 679 2842 735
rect 2898 679 2922 735
rect 2978 679 2984 735
rect 2836 642 2984 679
rect 54 433 82 485
rect 134 433 146 485
rect 198 433 231 485
rect 54 410 231 433
rect -805 378 -746 386
rect -805 322 -804 378
rect -748 322 -746 378
rect -805 298 -746 322
rect -805 242 -804 298
rect -748 242 -746 298
rect -805 234 -746 242
<< via2 >>
rect 2842 679 2898 735
rect 2922 679 2978 735
rect -804 322 -748 378
rect -804 242 -748 298
<< metal3 >>
rect 2828 735 2992 784
rect 2828 679 2842 735
rect 2898 679 2922 735
rect 2978 679 2992 735
rect 2828 564 2992 679
rect 2828 550 4095 564
rect 2828 486 4015 550
rect 4079 486 4095 550
rect 2828 470 4095 486
rect 2828 406 4015 470
rect 4079 406 4095 470
rect -1123 380 -738 395
rect 2828 391 4095 406
rect 2828 390 2992 391
rect -1123 316 -1078 380
rect -1014 378 -738 380
rect -1014 322 -804 378
rect -748 322 -738 378
rect -1014 316 -738 322
rect -1123 300 -738 316
rect -1123 236 -1078 300
rect -1014 298 -738 300
rect -1014 242 -804 298
rect -748 242 -738 298
rect -1014 236 -738 242
rect -1123 223 -738 236
<< via3 >>
rect 4015 486 4079 550
rect 4015 406 4079 470
rect -1078 316 -1014 380
rect -1078 236 -1014 300
<< metal4 >>
rect 3898 550 4098 566
rect 3898 486 4015 550
rect 4079 486 4098 550
rect 3898 470 4098 486
rect 3898 406 4015 470
rect 4079 406 4098 470
rect -1123 394 -968 395
rect -1952 380 -968 394
rect -1952 316 -1078 380
rect -1014 316 -968 380
rect -1952 300 -968 316
rect -1952 236 -1078 300
rect -1014 236 -968 300
rect -1952 231 -968 236
rect -1952 166 -976 231
rect -1952 -5924 -1704 166
rect 3898 -668 4098 406
rect -1784 -5930 -1704 -5924
use T_Gate  T_Gate_0
timestamp 1667803582
transform -1 0 -358 0 -1 2004
box -2642 0 541 1919
use T_Gate  T_Gate_1
timestamp 1667803582
transform 1 0 2642 0 1 0
box -2642 0 541 1919
use sky130_fd_pr__cap_mim_m3_1_MJDHVK  sky130_fd_pr__cap_mim_m3_1_MJDHVK_0
timestamp 1667803582
transform -1 0 1149 0 1 -3033
box -2950 -2900 2949 2900
use sky130_fd_pr__nfet_01v8_H73VBR  sky130_fd_pr__nfet_01v8_H73VBR_0
timestamp 1667803582
transform 1 0 200 0 1 2136
box -349 -450 349 450
<< labels >>
flabel metal2 s 579 2304 579 2304 0 FreeSans 2000 0 0 0 VGND
port 1 nsew
flabel metal1 s 488 1990 488 1990 0 FreeSans 2000 0 0 0 PH2
port 2 nsew
flabel metal3 s 3702 446 3702 446 0 FreeSans 2000 0 0 0 VOUT
port 3 nsew
<< end >>
