magic
tech sky130B
magscale 1 2
timestamp 1667803582
<< pwell >>
rect -415 1306 3823 1603
rect -415 -256 -109 1306
rect 3517 -256 3823 1306
rect -415 -553 3823 -256
<< psubdiff >>
rect -389 1573 3797 1577
rect -389 1335 375 1573
rect 3469 1335 3797 1573
rect -389 1332 3797 1335
rect -389 1028 -135 1332
rect -389 -26 -381 1028
rect -143 -26 -135 1028
rect 3543 1014 3797 1332
rect -389 -282 -135 -26
rect 3543 -40 3551 1014
rect 3789 -40 3797 1014
rect 3543 -282 3797 -40
rect -389 -286 3797 -282
rect -389 -524 33 -286
rect 3127 -524 3797 -286
rect -389 -527 3797 -524
<< psubdiffcont >>
rect 375 1335 3469 1573
rect -381 -26 -143 1028
rect 3551 -40 3789 1014
rect 33 -524 3127 -286
<< poly >>
rect 216 1144 3002 1158
rect 216 1110 250 1144
rect 284 1110 318 1144
rect 352 1110 386 1144
rect 420 1110 454 1144
rect 488 1110 522 1144
rect 556 1110 590 1144
rect 624 1110 658 1144
rect 692 1110 726 1144
rect 760 1110 794 1144
rect 828 1110 862 1144
rect 896 1110 930 1144
rect 964 1110 998 1144
rect 1032 1110 1066 1144
rect 1100 1110 1134 1144
rect 1168 1110 1202 1144
rect 1236 1110 1270 1144
rect 1304 1110 1338 1144
rect 1372 1110 1406 1144
rect 1440 1110 1474 1144
rect 1508 1110 1542 1144
rect 1576 1110 1610 1144
rect 1644 1110 1678 1144
rect 1712 1110 1746 1144
rect 1780 1110 1814 1144
rect 1848 1110 1882 1144
rect 1916 1110 1950 1144
rect 1984 1110 2018 1144
rect 2052 1110 2086 1144
rect 2120 1110 2154 1144
rect 2188 1110 2222 1144
rect 2256 1110 2290 1144
rect 2324 1110 2358 1144
rect 2392 1110 2426 1144
rect 2460 1110 2494 1144
rect 2528 1110 2562 1144
rect 2596 1110 2630 1144
rect 2664 1110 2698 1144
rect 2732 1110 2766 1144
rect 2800 1110 2834 1144
rect 2868 1110 2902 1144
rect 2936 1110 3002 1144
rect 216 1094 3002 1110
rect 216 1052 316 1094
rect 374 1052 474 1094
rect 848 1052 948 1094
rect 1006 1052 1106 1094
rect 1480 1052 1580 1094
rect 1638 1052 1738 1094
rect 2112 1052 2212 1094
rect 2270 1052 2370 1094
rect 2744 1052 2844 1094
rect 2902 1052 3002 1094
rect 58 -42 158 0
rect 532 -42 632 0
rect 690 -42 790 0
rect 1164 -42 1264 0
rect 1322 -42 1422 0
rect 1796 -42 1896 0
rect 1954 -42 2054 0
rect 2428 -42 2528 0
rect 2586 -42 2686 0
rect 3060 -42 3160 0
rect 58 -56 3160 -42
rect 58 -90 89 -56
rect 123 -90 157 -56
rect 191 -90 225 -56
rect 259 -90 293 -56
rect 327 -90 361 -56
rect 395 -90 429 -56
rect 463 -90 497 -56
rect 531 -90 565 -56
rect 599 -90 633 -56
rect 667 -90 701 -56
rect 735 -90 769 -56
rect 803 -90 837 -56
rect 871 -90 905 -56
rect 939 -90 973 -56
rect 1007 -90 1041 -56
rect 1075 -90 1109 -56
rect 1143 -90 1177 -56
rect 1211 -90 1245 -56
rect 1279 -90 1313 -56
rect 1347 -90 1381 -56
rect 1415 -90 1449 -56
rect 1483 -90 1517 -56
rect 1551 -90 1585 -56
rect 1619 -90 1653 -56
rect 1687 -90 1721 -56
rect 1755 -90 1789 -56
rect 1823 -90 1857 -56
rect 1891 -90 1925 -56
rect 1959 -90 1993 -56
rect 2027 -90 2061 -56
rect 2095 -90 2129 -56
rect 2163 -90 2197 -56
rect 2231 -90 2265 -56
rect 2299 -90 2333 -56
rect 2367 -90 2401 -56
rect 2435 -90 2469 -56
rect 2503 -90 2537 -56
rect 2571 -90 2605 -56
rect 2639 -90 2673 -56
rect 2707 -90 2741 -56
rect 2775 -90 2809 -56
rect 2843 -90 2877 -56
rect 2911 -90 2945 -56
rect 2979 -90 3013 -56
rect 3047 -90 3081 -56
rect 3115 -90 3160 -56
rect 58 -106 3160 -90
<< polycont >>
rect 250 1110 284 1144
rect 318 1110 352 1144
rect 386 1110 420 1144
rect 454 1110 488 1144
rect 522 1110 556 1144
rect 590 1110 624 1144
rect 658 1110 692 1144
rect 726 1110 760 1144
rect 794 1110 828 1144
rect 862 1110 896 1144
rect 930 1110 964 1144
rect 998 1110 1032 1144
rect 1066 1110 1100 1144
rect 1134 1110 1168 1144
rect 1202 1110 1236 1144
rect 1270 1110 1304 1144
rect 1338 1110 1372 1144
rect 1406 1110 1440 1144
rect 1474 1110 1508 1144
rect 1542 1110 1576 1144
rect 1610 1110 1644 1144
rect 1678 1110 1712 1144
rect 1746 1110 1780 1144
rect 1814 1110 1848 1144
rect 1882 1110 1916 1144
rect 1950 1110 1984 1144
rect 2018 1110 2052 1144
rect 2086 1110 2120 1144
rect 2154 1110 2188 1144
rect 2222 1110 2256 1144
rect 2290 1110 2324 1144
rect 2358 1110 2392 1144
rect 2426 1110 2460 1144
rect 2494 1110 2528 1144
rect 2562 1110 2596 1144
rect 2630 1110 2664 1144
rect 2698 1110 2732 1144
rect 2766 1110 2800 1144
rect 2834 1110 2868 1144
rect 2902 1110 2936 1144
rect 89 -90 123 -56
rect 157 -90 191 -56
rect 225 -90 259 -56
rect 293 -90 327 -56
rect 361 -90 395 -56
rect 429 -90 463 -56
rect 497 -90 531 -56
rect 565 -90 599 -56
rect 633 -90 667 -56
rect 701 -90 735 -56
rect 769 -90 803 -56
rect 837 -90 871 -56
rect 905 -90 939 -56
rect 973 -90 1007 -56
rect 1041 -90 1075 -56
rect 1109 -90 1143 -56
rect 1177 -90 1211 -56
rect 1245 -90 1279 -56
rect 1313 -90 1347 -56
rect 1381 -90 1415 -56
rect 1449 -90 1483 -56
rect 1517 -90 1551 -56
rect 1585 -90 1619 -56
rect 1653 -90 1687 -56
rect 1721 -90 1755 -56
rect 1789 -90 1823 -56
rect 1857 -90 1891 -56
rect 1925 -90 1959 -56
rect 1993 -90 2027 -56
rect 2061 -90 2095 -56
rect 2129 -90 2163 -56
rect 2197 -90 2231 -56
rect 2265 -90 2299 -56
rect 2333 -90 2367 -56
rect 2401 -90 2435 -56
rect 2469 -90 2503 -56
rect 2537 -90 2571 -56
rect 2605 -90 2639 -56
rect 2673 -90 2707 -56
rect 2741 -90 2775 -56
rect 2809 -90 2843 -56
rect 2877 -90 2911 -56
rect 2945 -90 2979 -56
rect 3013 -90 3047 -56
rect 3081 -90 3115 -56
<< locali >>
rect -389 1573 3797 1577
rect -389 1335 375 1573
rect 3469 1335 3797 1573
rect -389 1332 3797 1335
rect -389 1028 -135 1332
rect 216 1144 3002 1158
rect 216 1110 244 1144
rect 284 1110 316 1144
rect 352 1110 386 1144
rect 422 1110 454 1144
rect 494 1110 522 1144
rect 566 1110 590 1144
rect 638 1110 658 1144
rect 710 1110 726 1144
rect 782 1110 794 1144
rect 854 1110 862 1144
rect 926 1110 930 1144
rect 1032 1110 1036 1144
rect 1100 1110 1108 1144
rect 1168 1110 1180 1144
rect 1236 1110 1252 1144
rect 1304 1110 1324 1144
rect 1372 1110 1396 1144
rect 1440 1110 1468 1144
rect 1508 1110 1540 1144
rect 1576 1110 1610 1144
rect 1646 1110 1678 1144
rect 1718 1110 1746 1144
rect 1790 1110 1814 1144
rect 1862 1110 1882 1144
rect 1934 1110 1950 1144
rect 2006 1110 2018 1144
rect 2078 1110 2086 1144
rect 2150 1110 2154 1144
rect 2256 1110 2260 1144
rect 2324 1110 2332 1144
rect 2392 1110 2404 1144
rect 2460 1110 2476 1144
rect 2528 1110 2548 1144
rect 2596 1110 2620 1144
rect 2664 1110 2692 1144
rect 2732 1110 2764 1144
rect 2800 1110 2834 1144
rect 2870 1110 2902 1144
rect 2942 1110 3002 1144
rect 216 1094 3002 1110
rect -389 -26 -381 1028
rect -143 -26 -135 1028
rect -389 -282 -135 -26
rect 3543 1014 3797 1332
rect 3543 -40 3551 1014
rect 3789 -40 3797 1014
rect 58 -56 3160 -42
rect 58 -90 89 -56
rect 143 -90 157 -56
rect 215 -90 225 -56
rect 287 -90 293 -56
rect 359 -90 361 -56
rect 395 -90 397 -56
rect 463 -90 469 -56
rect 531 -90 541 -56
rect 599 -90 613 -56
rect 667 -90 685 -56
rect 735 -90 757 -56
rect 803 -90 829 -56
rect 871 -90 901 -56
rect 939 -90 973 -56
rect 1007 -90 1041 -56
rect 1079 -90 1109 -56
rect 1151 -90 1177 -56
rect 1223 -90 1245 -56
rect 1295 -90 1313 -56
rect 1367 -90 1381 -56
rect 1439 -90 1449 -56
rect 1511 -90 1517 -56
rect 1583 -90 1585 -56
rect 1619 -90 1621 -56
rect 1687 -90 1693 -56
rect 1755 -90 1765 -56
rect 1823 -90 1837 -56
rect 1891 -90 1909 -56
rect 1959 -90 1981 -56
rect 2027 -90 2053 -56
rect 2095 -90 2125 -56
rect 2163 -90 2197 -56
rect 2231 -90 2265 -56
rect 2303 -90 2333 -56
rect 2375 -90 2401 -56
rect 2447 -90 2469 -56
rect 2519 -90 2537 -56
rect 2591 -90 2605 -56
rect 2663 -90 2673 -56
rect 2735 -90 2741 -56
rect 2807 -90 2809 -56
rect 2843 -90 2845 -56
rect 2911 -90 2917 -56
rect 2979 -90 2989 -56
rect 3047 -90 3061 -56
rect 3115 -90 3160 -56
rect 58 -106 3160 -90
rect 3543 -282 3797 -40
rect -389 -286 3797 -282
rect -389 -524 33 -286
rect 3127 -524 3797 -286
rect -389 -527 3797 -524
<< viali >>
rect 244 1110 250 1144
rect 250 1110 278 1144
rect 316 1110 318 1144
rect 318 1110 350 1144
rect 388 1110 420 1144
rect 420 1110 422 1144
rect 460 1110 488 1144
rect 488 1110 494 1144
rect 532 1110 556 1144
rect 556 1110 566 1144
rect 604 1110 624 1144
rect 624 1110 638 1144
rect 676 1110 692 1144
rect 692 1110 710 1144
rect 748 1110 760 1144
rect 760 1110 782 1144
rect 820 1110 828 1144
rect 828 1110 854 1144
rect 892 1110 896 1144
rect 896 1110 926 1144
rect 964 1110 998 1144
rect 1036 1110 1066 1144
rect 1066 1110 1070 1144
rect 1108 1110 1134 1144
rect 1134 1110 1142 1144
rect 1180 1110 1202 1144
rect 1202 1110 1214 1144
rect 1252 1110 1270 1144
rect 1270 1110 1286 1144
rect 1324 1110 1338 1144
rect 1338 1110 1358 1144
rect 1396 1110 1406 1144
rect 1406 1110 1430 1144
rect 1468 1110 1474 1144
rect 1474 1110 1502 1144
rect 1540 1110 1542 1144
rect 1542 1110 1574 1144
rect 1612 1110 1644 1144
rect 1644 1110 1646 1144
rect 1684 1110 1712 1144
rect 1712 1110 1718 1144
rect 1756 1110 1780 1144
rect 1780 1110 1790 1144
rect 1828 1110 1848 1144
rect 1848 1110 1862 1144
rect 1900 1110 1916 1144
rect 1916 1110 1934 1144
rect 1972 1110 1984 1144
rect 1984 1110 2006 1144
rect 2044 1110 2052 1144
rect 2052 1110 2078 1144
rect 2116 1110 2120 1144
rect 2120 1110 2150 1144
rect 2188 1110 2222 1144
rect 2260 1110 2290 1144
rect 2290 1110 2294 1144
rect 2332 1110 2358 1144
rect 2358 1110 2366 1144
rect 2404 1110 2426 1144
rect 2426 1110 2438 1144
rect 2476 1110 2494 1144
rect 2494 1110 2510 1144
rect 2548 1110 2562 1144
rect 2562 1110 2582 1144
rect 2620 1110 2630 1144
rect 2630 1110 2654 1144
rect 2692 1110 2698 1144
rect 2698 1110 2726 1144
rect 2764 1110 2766 1144
rect 2766 1110 2798 1144
rect 2836 1110 2868 1144
rect 2868 1110 2870 1144
rect 2908 1110 2936 1144
rect 2936 1110 2942 1144
rect 109 -90 123 -56
rect 123 -90 143 -56
rect 181 -90 191 -56
rect 191 -90 215 -56
rect 253 -90 259 -56
rect 259 -90 287 -56
rect 325 -90 327 -56
rect 327 -90 359 -56
rect 397 -90 429 -56
rect 429 -90 431 -56
rect 469 -90 497 -56
rect 497 -90 503 -56
rect 541 -90 565 -56
rect 565 -90 575 -56
rect 613 -90 633 -56
rect 633 -90 647 -56
rect 685 -90 701 -56
rect 701 -90 719 -56
rect 757 -90 769 -56
rect 769 -90 791 -56
rect 829 -90 837 -56
rect 837 -90 863 -56
rect 901 -90 905 -56
rect 905 -90 935 -56
rect 973 -90 1007 -56
rect 1045 -90 1075 -56
rect 1075 -90 1079 -56
rect 1117 -90 1143 -56
rect 1143 -90 1151 -56
rect 1189 -90 1211 -56
rect 1211 -90 1223 -56
rect 1261 -90 1279 -56
rect 1279 -90 1295 -56
rect 1333 -90 1347 -56
rect 1347 -90 1367 -56
rect 1405 -90 1415 -56
rect 1415 -90 1439 -56
rect 1477 -90 1483 -56
rect 1483 -90 1511 -56
rect 1549 -90 1551 -56
rect 1551 -90 1583 -56
rect 1621 -90 1653 -56
rect 1653 -90 1655 -56
rect 1693 -90 1721 -56
rect 1721 -90 1727 -56
rect 1765 -90 1789 -56
rect 1789 -90 1799 -56
rect 1837 -90 1857 -56
rect 1857 -90 1871 -56
rect 1909 -90 1925 -56
rect 1925 -90 1943 -56
rect 1981 -90 1993 -56
rect 1993 -90 2015 -56
rect 2053 -90 2061 -56
rect 2061 -90 2087 -56
rect 2125 -90 2129 -56
rect 2129 -90 2159 -56
rect 2197 -90 2231 -56
rect 2269 -90 2299 -56
rect 2299 -90 2303 -56
rect 2341 -90 2367 -56
rect 2367 -90 2375 -56
rect 2413 -90 2435 -56
rect 2435 -90 2447 -56
rect 2485 -90 2503 -56
rect 2503 -90 2519 -56
rect 2557 -90 2571 -56
rect 2571 -90 2591 -56
rect 2629 -90 2639 -56
rect 2639 -90 2663 -56
rect 2701 -90 2707 -56
rect 2707 -90 2735 -56
rect 2773 -90 2775 -56
rect 2775 -90 2807 -56
rect 2845 -90 2877 -56
rect 2877 -90 2879 -56
rect 2917 -90 2945 -56
rect 2945 -90 2951 -56
rect 2989 -90 3013 -56
rect 3013 -90 3023 -56
rect 3061 -90 3081 -56
rect 3081 -90 3095 -56
<< metal1 >>
rect 216 1144 3002 1158
rect 216 1110 244 1144
rect 278 1110 316 1144
rect 350 1110 388 1144
rect 422 1110 460 1144
rect 494 1110 532 1144
rect 566 1110 604 1144
rect 638 1110 676 1144
rect 710 1110 748 1144
rect 782 1110 820 1144
rect 854 1110 892 1144
rect 926 1110 964 1144
rect 998 1110 1036 1144
rect 1070 1110 1108 1144
rect 1142 1110 1180 1144
rect 1214 1110 1252 1144
rect 1286 1110 1324 1144
rect 1358 1110 1396 1144
rect 1430 1110 1468 1144
rect 1502 1110 1540 1144
rect 1574 1110 1612 1144
rect 1646 1110 1684 1144
rect 1718 1110 1756 1144
rect 1790 1110 1828 1144
rect 1862 1110 1900 1144
rect 1934 1110 1972 1144
rect 2006 1110 2044 1144
rect 2078 1110 2116 1144
rect 2150 1110 2188 1144
rect 2222 1110 2260 1144
rect 2294 1110 2332 1144
rect 2366 1110 2404 1144
rect 2438 1110 2476 1144
rect 2510 1110 2548 1144
rect 2582 1110 2620 1144
rect 2654 1110 2692 1144
rect 2726 1110 2764 1144
rect 2798 1110 2836 1144
rect 2870 1110 2908 1144
rect 2942 1110 3002 1144
rect 216 1094 3002 1110
rect 313 928 377 959
rect 313 876 319 928
rect 371 876 377 928
rect 313 846 377 876
rect 945 928 1009 959
rect 945 876 951 928
rect 1003 876 1009 928
rect 945 846 1009 876
rect 1577 928 1641 959
rect 1577 876 1583 928
rect 1635 876 1641 928
rect 1577 846 1641 876
rect 2209 928 2273 959
rect 2209 876 2215 928
rect 2267 876 2273 928
rect 2209 846 2273 876
rect 2841 928 2905 959
rect 2841 876 2847 928
rect 2899 876 2905 928
rect 2841 846 2905 876
rect 158 585 216 619
rect 158 533 161 585
rect 213 533 216 585
rect 158 503 216 533
rect 474 585 532 619
rect 474 533 477 585
rect 529 533 532 585
rect 474 503 532 533
rect 790 585 848 619
rect 790 533 793 585
rect 845 533 848 585
rect 790 503 848 533
rect 1106 585 1164 619
rect 1106 533 1109 585
rect 1161 533 1164 585
rect 1106 503 1164 533
rect 1422 585 1480 619
rect 1422 533 1425 585
rect 1477 533 1480 585
rect 1422 503 1480 533
rect 1738 585 1796 619
rect 1738 533 1741 585
rect 1793 533 1796 585
rect 1738 503 1796 533
rect 2054 585 2112 619
rect 2054 533 2057 585
rect 2109 533 2112 585
rect 2054 503 2112 533
rect 2370 585 2428 619
rect 2370 533 2373 585
rect 2425 533 2428 585
rect 2370 503 2428 533
rect 2686 585 2744 619
rect 2686 533 2689 585
rect 2741 533 2744 585
rect 2686 503 2744 533
rect 3002 585 3060 619
rect 3002 533 3005 585
rect 3057 533 3060 585
rect 3002 503 3060 533
rect -3 156 61 188
rect -3 104 3 156
rect 55 104 61 156
rect -3 74 61 104
rect 629 156 693 188
rect 629 104 635 156
rect 687 104 693 156
rect 629 74 693 104
rect 1261 156 1325 188
rect 1261 104 1267 156
rect 1319 104 1325 156
rect 1261 74 1325 104
rect 1893 156 1957 188
rect 1893 104 1899 156
rect 1951 104 1957 156
rect 1893 74 1957 104
rect 2525 156 2589 188
rect 2525 104 2531 156
rect 2583 104 2589 156
rect 2525 74 2589 104
rect 3157 156 3221 188
rect 3157 104 3163 156
rect 3215 104 3221 156
rect 3157 74 3221 104
rect 58 -56 3160 -42
rect 58 -90 109 -56
rect 143 -90 181 -56
rect 215 -90 253 -56
rect 287 -90 325 -56
rect 359 -90 397 -56
rect 431 -90 469 -56
rect 503 -90 541 -56
rect 575 -90 613 -56
rect 647 -90 685 -56
rect 719 -90 757 -56
rect 791 -90 829 -56
rect 863 -90 901 -56
rect 935 -90 973 -56
rect 1007 -90 1045 -56
rect 1079 -90 1117 -56
rect 1151 -90 1189 -56
rect 1223 -90 1261 -56
rect 1295 -90 1333 -56
rect 1367 -90 1405 -56
rect 1439 -90 1477 -56
rect 1511 -90 1549 -56
rect 1583 -90 1621 -56
rect 1655 -90 1693 -56
rect 1727 -90 1765 -56
rect 1799 -90 1837 -56
rect 1871 -90 1909 -56
rect 1943 -90 1981 -56
rect 2015 -90 2053 -56
rect 2087 -90 2125 -56
rect 2159 -90 2197 -56
rect 2231 -90 2269 -56
rect 2303 -90 2341 -56
rect 2375 -90 2413 -56
rect 2447 -90 2485 -56
rect 2519 -90 2557 -56
rect 2591 -90 2629 -56
rect 2663 -90 2701 -56
rect 2735 -90 2773 -56
rect 2807 -90 2845 -56
rect 2879 -90 2917 -56
rect 2951 -90 2989 -56
rect 3023 -90 3061 -56
rect 3095 -90 3160 -56
rect 58 -106 3160 -90
<< via1 >>
rect 319 876 371 928
rect 951 876 1003 928
rect 1583 876 1635 928
rect 2215 876 2267 928
rect 2847 876 2899 928
rect 161 533 213 585
rect 477 533 529 585
rect 793 533 845 585
rect 1109 533 1161 585
rect 1425 533 1477 585
rect 1741 533 1793 585
rect 2057 533 2109 585
rect 2373 533 2425 585
rect 2689 533 2741 585
rect 3005 533 3057 585
rect 3 104 55 156
rect 635 104 687 156
rect 1267 104 1319 156
rect 1899 104 1951 156
rect 2531 104 2583 156
rect 3163 104 3215 156
<< metal2 >>
rect 0 928 3218 962
rect 0 876 319 928
rect 371 876 951 928
rect 1003 876 1583 928
rect 1635 876 2215 928
rect 2267 876 2847 928
rect 2899 876 3218 928
rect 0 846 3218 876
rect 0 585 3218 619
rect 0 533 161 585
rect 213 533 477 585
rect 529 533 793 585
rect 845 533 1109 585
rect 1161 533 1425 585
rect 1477 533 1741 585
rect 1793 533 2057 585
rect 2109 533 2373 585
rect 2425 533 2689 585
rect 2741 533 3005 585
rect 3057 533 3218 585
rect 0 503 3218 533
rect 0 156 3218 190
rect 0 104 3 156
rect 55 104 635 156
rect 687 104 1267 156
rect 1319 104 1899 156
rect 1951 104 2531 156
rect 2583 104 3163 156
rect 3215 104 3218 156
rect 0 74 3218 104
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_0
timestamp 1667803582
transform 1 0 3110 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_1
timestamp 1667803582
transform 1 0 2952 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_2
timestamp 1667803582
transform 1 0 2636 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_3
timestamp 1667803582
transform 1 0 2794 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_4
timestamp 1667803582
transform 1 0 2320 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_5
timestamp 1667803582
transform 1 0 2478 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_6
timestamp 1667803582
transform 1 0 2004 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_7
timestamp 1667803582
transform 1 0 2162 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_8
timestamp 1667803582
transform 1 0 1846 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_9
timestamp 1667803582
transform 1 0 1530 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_10
timestamp 1667803582
transform 1 0 1688 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_11
timestamp 1667803582
transform 1 0 1214 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_12
timestamp 1667803582
transform 1 0 1372 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_13
timestamp 1667803582
transform 1 0 1056 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_14
timestamp 1667803582
transform 1 0 740 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_15
timestamp 1667803582
transform 1 0 898 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_16
timestamp 1667803582
transform 1 0 424 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_17
timestamp 1667803582
transform 1 0 582 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_18
timestamp 1667803582
transform 1 0 108 0 1 526
box -134 -526 134 526
use sky130_fd_pr__nfet_01v8_6YBK2C  sky130_fd_pr__nfet_01v8_6YBK2C_19
timestamp 1667803582
transform 1 0 266 0 1 526
box -134 -526 134 526
<< labels >>
flabel metal1 s 408 -95 408 -95 0 FreeSans 1250 0 0 0 G1
port 1 nsew
flabel metal1 s 482 1139 482 1139 0 FreeSans 1250 0 0 0 G2
port 2 nsew
flabel metal2 s 3106 898 3106 898 0 FreeSans 1250 0 0 0 D2
port 3 nsew
flabel metal2 s 3111 542 3111 542 0 FreeSans 1250 0 0 0 S
port 4 nsew
flabel metal2 s 3085 128 3085 128 0 FreeSans 1250 0 0 0 D1
port 5 nsew
<< end >>
